//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[6][1]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Mon Jul  7 22:56:01 2025
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_6__1_ -----
module sb_6__1_(pReset,
                prog_clk,
                chany_top_in,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_,
                chany_bottom_in,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_2_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_3_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_4_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_5_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_6_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_7_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_8_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_9_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_10_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_11_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_12_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_13_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_14_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_15_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_16_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_17_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_18_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_19_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_20_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_21_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_22_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_23_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_24_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_25_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_26_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_27_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_28_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_29_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_30_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_31_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_32_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_33_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_34_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_35_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:149] chany_top_in;
//----- INPUT PORTS -----
input [0:149] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:149] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_2_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_3_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_4_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_5_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_6_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_7_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_8_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_9_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_10_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_11_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_12_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_13_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_14_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_15_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_16_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_17_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_18_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_19_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_20_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_21_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_22_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_23_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_24_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_25_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_26_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_27_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_28_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_29_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_30_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_31_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_32_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_33_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_34_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_35_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:149] chany_top_out;
//----- OUTPUT PORTS -----
output [0:149] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:149] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:7] mux_2level_tapbuf_size10_0_sram;
wire [0:7] mux_2level_tapbuf_size10_0_sram_inv;
wire [0:0] mux_2level_tapbuf_size10_mem_0_ccff_tail;
wire [0:7] mux_2level_tapbuf_size11_0_sram;
wire [0:7] mux_2level_tapbuf_size11_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_1_sram;
wire [0:7] mux_2level_tapbuf_size11_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_2_sram;
wire [0:7] mux_2level_tapbuf_size11_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_3_sram;
wire [0:7] mux_2level_tapbuf_size11_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_4_sram;
wire [0:7] mux_2level_tapbuf_size11_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_5_sram;
wire [0:7] mux_2level_tapbuf_size11_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_6_sram;
wire [0:7] mux_2level_tapbuf_size11_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_7_sram;
wire [0:7] mux_2level_tapbuf_size11_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_8_sram;
wire [0:7] mux_2level_tapbuf_size11_8_sram_inv;
wire [0:0] mux_2level_tapbuf_size11_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_8_ccff_tail;
wire [0:7] mux_2level_tapbuf_size12_0_sram;
wire [0:7] mux_2level_tapbuf_size12_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_10_sram;
wire [0:7] mux_2level_tapbuf_size12_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_11_sram;
wire [0:7] mux_2level_tapbuf_size12_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_12_sram;
wire [0:7] mux_2level_tapbuf_size12_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_13_sram;
wire [0:7] mux_2level_tapbuf_size12_13_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_14_sram;
wire [0:7] mux_2level_tapbuf_size12_14_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_15_sram;
wire [0:7] mux_2level_tapbuf_size12_15_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_16_sram;
wire [0:7] mux_2level_tapbuf_size12_16_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_17_sram;
wire [0:7] mux_2level_tapbuf_size12_17_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_18_sram;
wire [0:7] mux_2level_tapbuf_size12_18_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_19_sram;
wire [0:7] mux_2level_tapbuf_size12_19_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_1_sram;
wire [0:7] mux_2level_tapbuf_size12_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_20_sram;
wire [0:7] mux_2level_tapbuf_size12_20_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_21_sram;
wire [0:7] mux_2level_tapbuf_size12_21_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_22_sram;
wire [0:7] mux_2level_tapbuf_size12_22_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_23_sram;
wire [0:7] mux_2level_tapbuf_size12_23_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_24_sram;
wire [0:7] mux_2level_tapbuf_size12_24_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_25_sram;
wire [0:7] mux_2level_tapbuf_size12_25_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_26_sram;
wire [0:7] mux_2level_tapbuf_size12_26_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_2_sram;
wire [0:7] mux_2level_tapbuf_size12_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_3_sram;
wire [0:7] mux_2level_tapbuf_size12_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_4_sram;
wire [0:7] mux_2level_tapbuf_size12_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_5_sram;
wire [0:7] mux_2level_tapbuf_size12_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_6_sram;
wire [0:7] mux_2level_tapbuf_size12_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_7_sram;
wire [0:7] mux_2level_tapbuf_size12_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_8_sram;
wire [0:7] mux_2level_tapbuf_size12_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_9_sram;
wire [0:7] mux_2level_tapbuf_size12_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size12_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_9_ccff_tail;
wire [0:1] mux_2level_tapbuf_size3_0_sram;
wire [0:1] mux_2level_tapbuf_size3_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_100_sram;
wire [0:1] mux_2level_tapbuf_size3_100_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_101_sram;
wire [0:1] mux_2level_tapbuf_size3_101_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_102_sram;
wire [0:1] mux_2level_tapbuf_size3_102_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_103_sram;
wire [0:1] mux_2level_tapbuf_size3_103_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_104_sram;
wire [0:1] mux_2level_tapbuf_size3_104_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_105_sram;
wire [0:1] mux_2level_tapbuf_size3_105_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_106_sram;
wire [0:1] mux_2level_tapbuf_size3_106_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_107_sram;
wire [0:1] mux_2level_tapbuf_size3_107_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_108_sram;
wire [0:1] mux_2level_tapbuf_size3_108_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_109_sram;
wire [0:1] mux_2level_tapbuf_size3_109_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_10_sram;
wire [0:1] mux_2level_tapbuf_size3_10_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_110_sram;
wire [0:1] mux_2level_tapbuf_size3_110_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_111_sram;
wire [0:1] mux_2level_tapbuf_size3_111_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_112_sram;
wire [0:1] mux_2level_tapbuf_size3_112_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_113_sram;
wire [0:1] mux_2level_tapbuf_size3_113_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_114_sram;
wire [0:1] mux_2level_tapbuf_size3_114_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_115_sram;
wire [0:1] mux_2level_tapbuf_size3_115_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_116_sram;
wire [0:1] mux_2level_tapbuf_size3_116_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_117_sram;
wire [0:1] mux_2level_tapbuf_size3_117_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_118_sram;
wire [0:1] mux_2level_tapbuf_size3_118_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_119_sram;
wire [0:1] mux_2level_tapbuf_size3_119_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_11_sram;
wire [0:1] mux_2level_tapbuf_size3_11_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_120_sram;
wire [0:1] mux_2level_tapbuf_size3_120_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_121_sram;
wire [0:1] mux_2level_tapbuf_size3_121_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_122_sram;
wire [0:1] mux_2level_tapbuf_size3_122_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_123_sram;
wire [0:1] mux_2level_tapbuf_size3_123_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_124_sram;
wire [0:1] mux_2level_tapbuf_size3_124_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_125_sram;
wire [0:1] mux_2level_tapbuf_size3_125_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_126_sram;
wire [0:1] mux_2level_tapbuf_size3_126_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_127_sram;
wire [0:1] mux_2level_tapbuf_size3_127_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_128_sram;
wire [0:1] mux_2level_tapbuf_size3_128_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_129_sram;
wire [0:1] mux_2level_tapbuf_size3_129_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_12_sram;
wire [0:1] mux_2level_tapbuf_size3_12_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_130_sram;
wire [0:1] mux_2level_tapbuf_size3_130_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_131_sram;
wire [0:1] mux_2level_tapbuf_size3_131_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_132_sram;
wire [0:1] mux_2level_tapbuf_size3_132_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_133_sram;
wire [0:1] mux_2level_tapbuf_size3_133_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_134_sram;
wire [0:1] mux_2level_tapbuf_size3_134_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_135_sram;
wire [0:1] mux_2level_tapbuf_size3_135_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_136_sram;
wire [0:1] mux_2level_tapbuf_size3_136_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_137_sram;
wire [0:1] mux_2level_tapbuf_size3_137_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_138_sram;
wire [0:1] mux_2level_tapbuf_size3_138_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_139_sram;
wire [0:1] mux_2level_tapbuf_size3_139_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_13_sram;
wire [0:1] mux_2level_tapbuf_size3_13_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_140_sram;
wire [0:1] mux_2level_tapbuf_size3_140_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_141_sram;
wire [0:1] mux_2level_tapbuf_size3_141_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_142_sram;
wire [0:1] mux_2level_tapbuf_size3_142_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_143_sram;
wire [0:1] mux_2level_tapbuf_size3_143_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_14_sram;
wire [0:1] mux_2level_tapbuf_size3_14_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_15_sram;
wire [0:1] mux_2level_tapbuf_size3_15_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_16_sram;
wire [0:1] mux_2level_tapbuf_size3_16_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_17_sram;
wire [0:1] mux_2level_tapbuf_size3_17_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_18_sram;
wire [0:1] mux_2level_tapbuf_size3_18_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_19_sram;
wire [0:1] mux_2level_tapbuf_size3_19_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_1_sram;
wire [0:1] mux_2level_tapbuf_size3_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_20_sram;
wire [0:1] mux_2level_tapbuf_size3_20_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_21_sram;
wire [0:1] mux_2level_tapbuf_size3_21_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_22_sram;
wire [0:1] mux_2level_tapbuf_size3_22_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_23_sram;
wire [0:1] mux_2level_tapbuf_size3_23_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_24_sram;
wire [0:1] mux_2level_tapbuf_size3_24_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_25_sram;
wire [0:1] mux_2level_tapbuf_size3_25_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_26_sram;
wire [0:1] mux_2level_tapbuf_size3_26_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_27_sram;
wire [0:1] mux_2level_tapbuf_size3_27_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_28_sram;
wire [0:1] mux_2level_tapbuf_size3_28_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_29_sram;
wire [0:1] mux_2level_tapbuf_size3_29_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_2_sram;
wire [0:1] mux_2level_tapbuf_size3_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_30_sram;
wire [0:1] mux_2level_tapbuf_size3_30_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_31_sram;
wire [0:1] mux_2level_tapbuf_size3_31_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_32_sram;
wire [0:1] mux_2level_tapbuf_size3_32_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_33_sram;
wire [0:1] mux_2level_tapbuf_size3_33_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_34_sram;
wire [0:1] mux_2level_tapbuf_size3_34_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_35_sram;
wire [0:1] mux_2level_tapbuf_size3_35_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_36_sram;
wire [0:1] mux_2level_tapbuf_size3_36_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_37_sram;
wire [0:1] mux_2level_tapbuf_size3_37_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_38_sram;
wire [0:1] mux_2level_tapbuf_size3_38_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_39_sram;
wire [0:1] mux_2level_tapbuf_size3_39_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_3_sram;
wire [0:1] mux_2level_tapbuf_size3_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_40_sram;
wire [0:1] mux_2level_tapbuf_size3_40_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_41_sram;
wire [0:1] mux_2level_tapbuf_size3_41_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_42_sram;
wire [0:1] mux_2level_tapbuf_size3_42_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_43_sram;
wire [0:1] mux_2level_tapbuf_size3_43_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_44_sram;
wire [0:1] mux_2level_tapbuf_size3_44_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_45_sram;
wire [0:1] mux_2level_tapbuf_size3_45_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_46_sram;
wire [0:1] mux_2level_tapbuf_size3_46_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_47_sram;
wire [0:1] mux_2level_tapbuf_size3_47_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_48_sram;
wire [0:1] mux_2level_tapbuf_size3_48_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_49_sram;
wire [0:1] mux_2level_tapbuf_size3_49_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_4_sram;
wire [0:1] mux_2level_tapbuf_size3_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_50_sram;
wire [0:1] mux_2level_tapbuf_size3_50_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_51_sram;
wire [0:1] mux_2level_tapbuf_size3_51_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_52_sram;
wire [0:1] mux_2level_tapbuf_size3_52_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_53_sram;
wire [0:1] mux_2level_tapbuf_size3_53_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_54_sram;
wire [0:1] mux_2level_tapbuf_size3_54_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_55_sram;
wire [0:1] mux_2level_tapbuf_size3_55_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_56_sram;
wire [0:1] mux_2level_tapbuf_size3_56_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_57_sram;
wire [0:1] mux_2level_tapbuf_size3_57_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_58_sram;
wire [0:1] mux_2level_tapbuf_size3_58_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_59_sram;
wire [0:1] mux_2level_tapbuf_size3_59_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_5_sram;
wire [0:1] mux_2level_tapbuf_size3_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_60_sram;
wire [0:1] mux_2level_tapbuf_size3_60_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_61_sram;
wire [0:1] mux_2level_tapbuf_size3_61_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_62_sram;
wire [0:1] mux_2level_tapbuf_size3_62_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_63_sram;
wire [0:1] mux_2level_tapbuf_size3_63_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_64_sram;
wire [0:1] mux_2level_tapbuf_size3_64_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_65_sram;
wire [0:1] mux_2level_tapbuf_size3_65_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_66_sram;
wire [0:1] mux_2level_tapbuf_size3_66_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_67_sram;
wire [0:1] mux_2level_tapbuf_size3_67_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_68_sram;
wire [0:1] mux_2level_tapbuf_size3_68_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_69_sram;
wire [0:1] mux_2level_tapbuf_size3_69_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_6_sram;
wire [0:1] mux_2level_tapbuf_size3_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_70_sram;
wire [0:1] mux_2level_tapbuf_size3_70_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_71_sram;
wire [0:1] mux_2level_tapbuf_size3_71_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_72_sram;
wire [0:1] mux_2level_tapbuf_size3_72_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_73_sram;
wire [0:1] mux_2level_tapbuf_size3_73_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_74_sram;
wire [0:1] mux_2level_tapbuf_size3_74_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_75_sram;
wire [0:1] mux_2level_tapbuf_size3_75_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_76_sram;
wire [0:1] mux_2level_tapbuf_size3_76_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_77_sram;
wire [0:1] mux_2level_tapbuf_size3_77_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_78_sram;
wire [0:1] mux_2level_tapbuf_size3_78_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_79_sram;
wire [0:1] mux_2level_tapbuf_size3_79_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_7_sram;
wire [0:1] mux_2level_tapbuf_size3_7_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_80_sram;
wire [0:1] mux_2level_tapbuf_size3_80_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_81_sram;
wire [0:1] mux_2level_tapbuf_size3_81_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_82_sram;
wire [0:1] mux_2level_tapbuf_size3_82_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_83_sram;
wire [0:1] mux_2level_tapbuf_size3_83_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_84_sram;
wire [0:1] mux_2level_tapbuf_size3_84_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_85_sram;
wire [0:1] mux_2level_tapbuf_size3_85_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_86_sram;
wire [0:1] mux_2level_tapbuf_size3_86_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_87_sram;
wire [0:1] mux_2level_tapbuf_size3_87_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_88_sram;
wire [0:1] mux_2level_tapbuf_size3_88_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_89_sram;
wire [0:1] mux_2level_tapbuf_size3_89_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_8_sram;
wire [0:1] mux_2level_tapbuf_size3_8_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_90_sram;
wire [0:1] mux_2level_tapbuf_size3_90_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_91_sram;
wire [0:1] mux_2level_tapbuf_size3_91_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_92_sram;
wire [0:1] mux_2level_tapbuf_size3_92_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_93_sram;
wire [0:1] mux_2level_tapbuf_size3_93_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_94_sram;
wire [0:1] mux_2level_tapbuf_size3_94_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_95_sram;
wire [0:1] mux_2level_tapbuf_size3_95_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_96_sram;
wire [0:1] mux_2level_tapbuf_size3_96_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_97_sram;
wire [0:1] mux_2level_tapbuf_size3_97_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_98_sram;
wire [0:1] mux_2level_tapbuf_size3_98_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_99_sram;
wire [0:1] mux_2level_tapbuf_size3_99_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_9_sram;
wire [0:1] mux_2level_tapbuf_size3_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_100_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_101_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_102_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_103_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_104_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_105_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_106_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_107_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_108_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_109_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_110_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_111_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_112_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_113_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_114_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_115_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_116_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_117_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_118_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_119_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_120_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_121_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_122_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_123_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_124_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_125_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_126_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_127_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_128_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_129_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_130_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_131_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_132_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_133_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_134_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_135_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_136_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_137_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_138_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_139_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_140_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_141_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_142_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_143_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_79_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_80_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_81_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_82_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_83_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_84_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_85_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_86_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_87_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_88_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_89_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_90_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_91_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_92_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_93_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_94_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_95_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_96_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_97_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_98_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_99_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size4_0_sram;
wire [0:5] mux_2level_tapbuf_size4_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_1_sram;
wire [0:5] mux_2level_tapbuf_size4_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_2_sram;
wire [0:5] mux_2level_tapbuf_size4_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_3_sram;
wire [0:5] mux_2level_tapbuf_size4_3_sram_inv;
wire [0:0] mux_2level_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_3_ccff_tail;
wire [0:5] mux_2level_tapbuf_size5_0_sram;
wire [0:5] mux_2level_tapbuf_size5_0_sram_inv;
wire [0:0] mux_2level_tapbuf_size5_mem_0_ccff_tail;
wire [0:5] mux_2level_tapbuf_size6_0_sram;
wire [0:5] mux_2level_tapbuf_size6_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_1_sram;
wire [0:5] mux_2level_tapbuf_size6_1_sram_inv;
wire [0:0] mux_2level_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_1_ccff_tail;
wire [0:5] mux_2level_tapbuf_size7_0_sram;
wire [0:5] mux_2level_tapbuf_size7_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_10_sram;
wire [0:5] mux_2level_tapbuf_size7_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_11_sram;
wire [0:5] mux_2level_tapbuf_size7_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_12_sram;
wire [0:5] mux_2level_tapbuf_size7_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_13_sram;
wire [0:5] mux_2level_tapbuf_size7_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_14_sram;
wire [0:5] mux_2level_tapbuf_size7_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_15_sram;
wire [0:5] mux_2level_tapbuf_size7_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_16_sram;
wire [0:5] mux_2level_tapbuf_size7_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_17_sram;
wire [0:5] mux_2level_tapbuf_size7_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_18_sram;
wire [0:5] mux_2level_tapbuf_size7_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_19_sram;
wire [0:5] mux_2level_tapbuf_size7_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_1_sram;
wire [0:5] mux_2level_tapbuf_size7_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_20_sram;
wire [0:5] mux_2level_tapbuf_size7_20_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_21_sram;
wire [0:5] mux_2level_tapbuf_size7_21_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_22_sram;
wire [0:5] mux_2level_tapbuf_size7_22_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_23_sram;
wire [0:5] mux_2level_tapbuf_size7_23_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_24_sram;
wire [0:5] mux_2level_tapbuf_size7_24_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_25_sram;
wire [0:5] mux_2level_tapbuf_size7_25_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_26_sram;
wire [0:5] mux_2level_tapbuf_size7_26_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_27_sram;
wire [0:5] mux_2level_tapbuf_size7_27_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_28_sram;
wire [0:5] mux_2level_tapbuf_size7_28_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_29_sram;
wire [0:5] mux_2level_tapbuf_size7_29_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_2_sram;
wire [0:5] mux_2level_tapbuf_size7_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_30_sram;
wire [0:5] mux_2level_tapbuf_size7_30_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_31_sram;
wire [0:5] mux_2level_tapbuf_size7_31_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_32_sram;
wire [0:5] mux_2level_tapbuf_size7_32_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_33_sram;
wire [0:5] mux_2level_tapbuf_size7_33_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_34_sram;
wire [0:5] mux_2level_tapbuf_size7_34_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_3_sram;
wire [0:5] mux_2level_tapbuf_size7_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_4_sram;
wire [0:5] mux_2level_tapbuf_size7_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_5_sram;
wire [0:5] mux_2level_tapbuf_size7_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_6_sram;
wire [0:5] mux_2level_tapbuf_size7_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_7_sram;
wire [0:5] mux_2level_tapbuf_size7_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_8_sram;
wire [0:5] mux_2level_tapbuf_size7_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_9_sram;
wire [0:5] mux_2level_tapbuf_size7_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_9_ccff_tail;
wire [0:7] mux_2level_tapbuf_size9_0_sram;
wire [0:7] mux_2level_tapbuf_size9_0_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[105] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[106] = chany_top_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[109] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[110] = chany_top_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[111] = chany_top_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[113] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[114] = chany_top_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[115] = chany_top_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[117] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[118] = chany_top_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[119] = chany_top_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[121] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[122] = chany_top_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[123] = chany_top_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[126] = chany_top_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[127] = chany_top_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[129] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[130] = chany_top_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[131] = chany_top_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[133] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[135] = chany_top_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[137] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[138] = chany_top_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[139] = chany_top_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[141] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[142] = chany_top_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[145] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[146] = chany_top_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[147] = chany_top_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[149] = chany_top_in[148];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[0] = right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_[0];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 14 -----
	assign chanx_right_out[149] = right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_[0];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 330 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 334 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 338 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 342 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[105] = chany_bottom_in[104];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[106] = chany_bottom_in[105];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[107] = chany_bottom_in[106];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[109] = chany_bottom_in[108];
// ----- Local connection due to Wire 419 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[110] = chany_bottom_in[109];
// ----- Local connection due to Wire 420 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[111] = chany_bottom_in[110];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[113] = chany_bottom_in[112];
// ----- Local connection due to Wire 423 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[114] = chany_bottom_in[113];
// ----- Local connection due to Wire 424 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[115] = chany_bottom_in[114];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[117] = chany_bottom_in[116];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[118] = chany_bottom_in[117];
// ----- Local connection due to Wire 428 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[119] = chany_bottom_in[118];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[121] = chany_bottom_in[120];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[122] = chany_bottom_in[121];
// ----- Local connection due to Wire 432 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[123] = chany_bottom_in[122];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[125] = chany_bottom_in[124];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[126] = chany_bottom_in[125];
// ----- Local connection due to Wire 436 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[127] = chany_bottom_in[126];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[129] = chany_bottom_in[128];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[130] = chany_bottom_in[129];
// ----- Local connection due to Wire 440 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[131] = chany_bottom_in[130];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[133] = chany_bottom_in[132];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[134] = chany_bottom_in[133];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[135] = chany_bottom_in[134];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[137] = chany_bottom_in[136];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[138] = chany_bottom_in[137];
// ----- Local connection due to Wire 448 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[139] = chany_bottom_in[138];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[141] = chany_bottom_in[140];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[142] = chany_bottom_in[141];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[143] = chany_bottom_in[142];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[145] = chany_bottom_in[144];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[146] = chany_bottom_in[145];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[147] = chany_bottom_in[146];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[149] = chany_bottom_in[148];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size7 mux_top_track_0 (
		.in({chanx_right_in[1], chanx_right_in[39], chanx_right_in[77], chanx_right_in[115], chany_bottom_in[0], chany_bottom_in[50], chany_bottom_in[101]}),
		.sram(mux_2level_tapbuf_size7_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_0_sram_inv[0:5]),
		.out(chany_top_out[0]));

	mux_2level_tapbuf_size7 mux_top_track_8 (
		.in({chanx_right_in[2], chanx_right_in[40], chanx_right_in[78], chanx_right_in[116], chany_bottom_in[1], chany_bottom_in[52], chany_bottom_in[102]}),
		.sram(mux_2level_tapbuf_size7_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_1_sram_inv[0:5]),
		.out(chany_top_out[4]));

	mux_2level_tapbuf_size7 mux_top_track_16 (
		.in({chanx_right_in[3], chanx_right_in[41], chanx_right_in[79], chanx_right_in[117], chany_bottom_in[2], chany_bottom_in[53], chany_bottom_in[104]}),
		.sram(mux_2level_tapbuf_size7_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_2_sram_inv[0:5]),
		.out(chany_top_out[8]));

	mux_2level_tapbuf_size7 mux_top_track_24 (
		.in({chanx_right_in[4], chanx_right_in[42], chanx_right_in[80], chanx_right_in[118], chany_bottom_in[4], chany_bottom_in[54], chany_bottom_in[105]}),
		.sram(mux_2level_tapbuf_size7_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_3_sram_inv[0:5]),
		.out(chany_top_out[12]));

	mux_2level_tapbuf_size7 mux_top_track_32 (
		.in({chanx_right_in[5], chanx_right_in[43], chanx_right_in[81], chanx_right_in[119], chany_bottom_in[5], chany_bottom_in[56], chany_bottom_in[106]}),
		.sram(mux_2level_tapbuf_size7_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_4_sram_inv[0:5]),
		.out(chany_top_out[16]));

	mux_2level_tapbuf_size7 mux_top_track_40 (
		.in({chanx_right_in[6], chanx_right_in[44], chanx_right_in[82], chanx_right_in[120], chany_bottom_in[6], chany_bottom_in[57], chany_bottom_in[108]}),
		.sram(mux_2level_tapbuf_size7_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_5_sram_inv[0:5]),
		.out(chany_top_out[20]));

	mux_2level_tapbuf_size7 mux_top_track_48 (
		.in({chanx_right_in[7], chanx_right_in[45], chanx_right_in[83], chanx_right_in[121], chany_bottom_in[8], chany_bottom_in[58], chany_bottom_in[109]}),
		.sram(mux_2level_tapbuf_size7_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_6_sram_inv[0:5]),
		.out(chany_top_out[24]));

	mux_2level_tapbuf_size7 mux_top_track_56 (
		.in({chanx_right_in[8], chanx_right_in[46], chanx_right_in[84], chanx_right_in[122], chany_bottom_in[9], chany_bottom_in[60], chany_bottom_in[110]}),
		.sram(mux_2level_tapbuf_size7_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_7_sram_inv[0:5]),
		.out(chany_top_out[28]));

	mux_2level_tapbuf_size7 mux_top_track_64 (
		.in({chanx_right_in[9], chanx_right_in[47], chanx_right_in[85], chanx_right_in[123], chany_bottom_in[10], chany_bottom_in[61], chany_bottom_in[112]}),
		.sram(mux_2level_tapbuf_size7_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_8_sram_inv[0:5]),
		.out(chany_top_out[32]));

	mux_2level_tapbuf_size7 mux_top_track_72 (
		.in({chanx_right_in[10], chanx_right_in[48], chanx_right_in[86], chanx_right_in[124], chany_bottom_in[12], chany_bottom_in[62], chany_bottom_in[113]}),
		.sram(mux_2level_tapbuf_size7_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_9_sram_inv[0:5]),
		.out(chany_top_out[36]));

	mux_2level_tapbuf_size7 mux_top_track_80 (
		.in({chanx_right_in[11], chanx_right_in[49], chanx_right_in[87], chanx_right_in[125], chany_bottom_in[13], chany_bottom_in[64], chany_bottom_in[114]}),
		.sram(mux_2level_tapbuf_size7_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_10_sram_inv[0:5]),
		.out(chany_top_out[40]));

	mux_2level_tapbuf_size7 mux_top_track_88 (
		.in({chanx_right_in[12], chanx_right_in[50], chanx_right_in[88], chanx_right_in[126], chany_bottom_in[14], chany_bottom_in[65], chany_bottom_in[116]}),
		.sram(mux_2level_tapbuf_size7_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_11_sram_inv[0:5]),
		.out(chany_top_out[44]));

	mux_2level_tapbuf_size7 mux_top_track_96 (
		.in({chanx_right_in[13], chanx_right_in[51], chanx_right_in[89], chanx_right_in[127], chany_bottom_in[16], chany_bottom_in[66], chany_bottom_in[117]}),
		.sram(mux_2level_tapbuf_size7_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_12_sram_inv[0:5]),
		.out(chany_top_out[48]));

	mux_2level_tapbuf_size7 mux_top_track_104 (
		.in({chanx_right_in[14], chanx_right_in[52], chanx_right_in[90], chanx_right_in[128], chany_bottom_in[17], chany_bottom_in[68], chany_bottom_in[118]}),
		.sram(mux_2level_tapbuf_size7_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_13_sram_inv[0:5]),
		.out(chany_top_out[52]));

	mux_2level_tapbuf_size7 mux_top_track_112 (
		.in({chanx_right_in[15], chanx_right_in[53], chanx_right_in[91], chanx_right_in[129], chany_bottom_in[18], chany_bottom_in[69], chany_bottom_in[120]}),
		.sram(mux_2level_tapbuf_size7_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_14_sram_inv[0:5]),
		.out(chany_top_out[56]));

	mux_2level_tapbuf_size7 mux_top_track_120 (
		.in({chanx_right_in[16], chanx_right_in[54], chanx_right_in[92], chanx_right_in[130], chany_bottom_in[20], chany_bottom_in[70], chany_bottom_in[121]}),
		.sram(mux_2level_tapbuf_size7_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_15_sram_inv[0:5]),
		.out(chany_top_out[60]));

	mux_2level_tapbuf_size7 mux_top_track_128 (
		.in({chanx_right_in[17], chanx_right_in[55], chanx_right_in[93], chanx_right_in[131], chany_bottom_in[21], chany_bottom_in[72], chany_bottom_in[122]}),
		.sram(mux_2level_tapbuf_size7_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_16_sram_inv[0:5]),
		.out(chany_top_out[64]));

	mux_2level_tapbuf_size7 mux_top_track_136 (
		.in({chanx_right_in[18], chanx_right_in[56], chanx_right_in[94], chanx_right_in[132], chany_bottom_in[22], chany_bottom_in[73], chany_bottom_in[124]}),
		.sram(mux_2level_tapbuf_size7_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_17_sram_inv[0:5]),
		.out(chany_top_out[68]));

	mux_2level_tapbuf_size7 mux_top_track_144 (
		.in({chanx_right_in[19], chanx_right_in[57], chanx_right_in[95], chanx_right_in[133], chany_bottom_in[24], chany_bottom_in[74], chany_bottom_in[125]}),
		.sram(mux_2level_tapbuf_size7_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_18_sram_inv[0:5]),
		.out(chany_top_out[72]));

	mux_2level_tapbuf_size7 mux_top_track_152 (
		.in({chanx_right_in[20], chanx_right_in[58], chanx_right_in[96], chanx_right_in[134], chany_bottom_in[25], chany_bottom_in[76], chany_bottom_in[126]}),
		.sram(mux_2level_tapbuf_size7_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_19_sram_inv[0:5]),
		.out(chany_top_out[76]));

	mux_2level_tapbuf_size7 mux_top_track_160 (
		.in({chanx_right_in[21], chanx_right_in[59], chanx_right_in[97], chanx_right_in[135], chany_bottom_in[26], chany_bottom_in[77], chany_bottom_in[128]}),
		.sram(mux_2level_tapbuf_size7_20_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_20_sram_inv[0:5]),
		.out(chany_top_out[80]));

	mux_2level_tapbuf_size7 mux_top_track_168 (
		.in({chanx_right_in[22], chanx_right_in[60], chanx_right_in[98], chanx_right_in[136], chany_bottom_in[28], chany_bottom_in[78], chany_bottom_in[129]}),
		.sram(mux_2level_tapbuf_size7_21_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_21_sram_inv[0:5]),
		.out(chany_top_out[84]));

	mux_2level_tapbuf_size7 mux_top_track_176 (
		.in({chanx_right_in[23], chanx_right_in[61], chanx_right_in[99], chanx_right_in[137], chany_bottom_in[29], chany_bottom_in[80], chany_bottom_in[130]}),
		.sram(mux_2level_tapbuf_size7_22_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_22_sram_inv[0:5]),
		.out(chany_top_out[88]));

	mux_2level_tapbuf_size7 mux_top_track_184 (
		.in({chanx_right_in[24], chanx_right_in[62], chanx_right_in[100], chanx_right_in[138], chany_bottom_in[30], chany_bottom_in[81], chany_bottom_in[132]}),
		.sram(mux_2level_tapbuf_size7_23_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_23_sram_inv[0:5]),
		.out(chany_top_out[92]));

	mux_2level_tapbuf_size7 mux_top_track_192 (
		.in({chanx_right_in[25], chanx_right_in[63], chanx_right_in[101], chanx_right_in[139], chany_bottom_in[32], chany_bottom_in[82], chany_bottom_in[133]}),
		.sram(mux_2level_tapbuf_size7_24_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_24_sram_inv[0:5]),
		.out(chany_top_out[96]));

	mux_2level_tapbuf_size7 mux_top_track_200 (
		.in({chanx_right_in[26], chanx_right_in[64], chanx_right_in[102], chanx_right_in[140], chany_bottom_in[33], chany_bottom_in[84], chany_bottom_in[134]}),
		.sram(mux_2level_tapbuf_size7_25_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_25_sram_inv[0:5]),
		.out(chany_top_out[100]));

	mux_2level_tapbuf_size7 mux_top_track_208 (
		.in({chanx_right_in[27], chanx_right_in[65], chanx_right_in[103], chanx_right_in[141], chany_bottom_in[34], chany_bottom_in[85], chany_bottom_in[136]}),
		.sram(mux_2level_tapbuf_size7_26_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_26_sram_inv[0:5]),
		.out(chany_top_out[104]));

	mux_2level_tapbuf_size7 mux_top_track_216 (
		.in({chanx_right_in[28], chanx_right_in[66], chanx_right_in[104], chanx_right_in[142], chany_bottom_in[36], chany_bottom_in[86], chany_bottom_in[137]}),
		.sram(mux_2level_tapbuf_size7_27_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_27_sram_inv[0:5]),
		.out(chany_top_out[108]));

	mux_2level_tapbuf_size7 mux_top_track_224 (
		.in({chanx_right_in[29], chanx_right_in[67], chanx_right_in[105], chanx_right_in[143], chany_bottom_in[37], chany_bottom_in[88], chany_bottom_in[138]}),
		.sram(mux_2level_tapbuf_size7_28_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_28_sram_inv[0:5]),
		.out(chany_top_out[112]));

	mux_2level_tapbuf_size7 mux_top_track_232 (
		.in({chanx_right_in[30], chanx_right_in[68], chanx_right_in[106], chanx_right_in[144], chany_bottom_in[38], chany_bottom_in[89], chany_bottom_in[140]}),
		.sram(mux_2level_tapbuf_size7_29_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_29_sram_inv[0:5]),
		.out(chany_top_out[116]));

	mux_2level_tapbuf_size7 mux_top_track_240 (
		.in({chanx_right_in[31], chanx_right_in[69], chanx_right_in[107], chanx_right_in[145], chany_bottom_in[40], chany_bottom_in[90], chany_bottom_in[141]}),
		.sram(mux_2level_tapbuf_size7_30_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_30_sram_inv[0:5]),
		.out(chany_top_out[120]));

	mux_2level_tapbuf_size7 mux_top_track_248 (
		.in({chanx_right_in[32], chanx_right_in[70], chanx_right_in[108], chanx_right_in[146], chany_bottom_in[41], chany_bottom_in[92], chany_bottom_in[142]}),
		.sram(mux_2level_tapbuf_size7_31_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_31_sram_inv[0:5]),
		.out(chany_top_out[124]));

	mux_2level_tapbuf_size7 mux_top_track_256 (
		.in({chanx_right_in[33], chanx_right_in[71], chanx_right_in[109], chanx_right_in[147], chany_bottom_in[42], chany_bottom_in[93], chany_bottom_in[144]}),
		.sram(mux_2level_tapbuf_size7_32_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_32_sram_inv[0:5]),
		.out(chany_top_out[128]));

	mux_2level_tapbuf_size7 mux_top_track_264 (
		.in({chanx_right_in[34], chanx_right_in[72], chanx_right_in[110], chanx_right_in[148], chany_bottom_in[44], chany_bottom_in[94], chany_bottom_in[145]}),
		.sram(mux_2level_tapbuf_size7_33_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_33_sram_inv[0:5]),
		.out(chany_top_out[132]));

	mux_2level_tapbuf_size7 mux_top_track_272 (
		.in({chanx_right_in[35], chanx_right_in[73], chanx_right_in[111], chanx_right_in[149], chany_bottom_in[45], chany_bottom_in[96], chany_bottom_in[146]}),
		.sram(mux_2level_tapbuf_size7_34_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_34_sram_inv[0:5]),
		.out(chany_top_out[136]));

	mux_2level_tapbuf_size7_mem mem_top_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_0_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_1_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_2_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_3_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_4_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_5_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_6_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_7_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_8_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_9_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_10_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_11_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_12_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_13_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_14_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_15_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_16_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_17_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_18_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_19_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_20_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_20_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_21_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_21_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_22_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_22_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_23_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_23_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_24_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_24_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_25_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_25_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_26_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_26_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_27_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_27_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_28_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_28_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_29_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_29_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_30_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_30_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_31_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_31_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_32_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_32_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_33_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_33_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_34_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_34_sram_inv[0:5]));

	mux_2level_tapbuf_size6 mux_top_track_280 (
		.in({chanx_right_in[36], chanx_right_in[74], chanx_right_in[112], chany_bottom_in[46], chany_bottom_in[97], chany_bottom_in[148]}),
		.sram(mux_2level_tapbuf_size6_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_0_sram_inv[0:5]),
		.out(chany_top_out[140]));

	mux_2level_tapbuf_size6 mux_top_track_296 (
		.in({chanx_right_in[0], chanx_right_in[38], chanx_right_in[76], chanx_right_in[114], chany_bottom_in[49], chany_bottom_in[100]}),
		.sram(mux_2level_tapbuf_size6_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_1_sram_inv[0:5]),
		.out(chany_top_out[148]));

	mux_2level_tapbuf_size6_mem mem_top_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_0_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_1_sram_inv[0:5]));

	mux_2level_tapbuf_size5 mux_top_track_288 (
		.in({chanx_right_in[37], chanx_right_in[75], chanx_right_in[113], chany_bottom_in[48], chany_bottom_in[98]}),
		.sram(mux_2level_tapbuf_size5_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_0_sram_inv[0:5]),
		.out(chany_top_out[144]));

	mux_2level_tapbuf_size5_mem mem_top_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_0_sram_inv[0:5]));

	mux_2level_tapbuf_size3 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[3], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_}),
		.sram(mux_2level_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_0_sram_inv[0:1]),
		.out(chanx_right_out[1]));

	mux_2level_tapbuf_size3 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[7], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_1_sram_inv[0:1]),
		.out(chanx_right_out[2]));

	mux_2level_tapbuf_size3 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[11], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_}),
		.sram(mux_2level_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_2_sram_inv[0:1]),
		.out(chanx_right_out[3]));

	mux_2level_tapbuf_size3 mux_right_track_8 (
		.in({chany_top_in[4], chany_top_in[15], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_}),
		.sram(mux_2level_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_3_sram_inv[0:1]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size3 mux_right_track_10 (
		.in({chany_top_in[5], chany_top_in[19], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_}),
		.sram(mux_2level_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_4_sram_inv[0:1]),
		.out(chanx_right_out[5]));

	mux_2level_tapbuf_size3 mux_right_track_12 (
		.in({chany_top_in[6], chany_top_in[23], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_5_sram_inv[0:1]),
		.out(chanx_right_out[6]));

	mux_2level_tapbuf_size3 mux_right_track_14 (
		.in({chany_top_in[8], chany_top_in[27], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_}),
		.sram(mux_2level_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_6_sram_inv[0:1]),
		.out(chanx_right_out[7]));

	mux_2level_tapbuf_size3 mux_right_track_16 (
		.in({chany_top_in[9], chany_top_in[31], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_7_sram_inv[0:1]),
		.out(chanx_right_out[8]));

	mux_2level_tapbuf_size3 mux_right_track_18 (
		.in({chany_top_in[10], chany_top_in[35], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_8_sram_inv[0:1]),
		.out(chanx_right_out[9]));

	mux_2level_tapbuf_size3 mux_right_track_20 (
		.in({chany_top_in[12], chany_top_in[39], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_}),
		.sram(mux_2level_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_9_sram_inv[0:1]),
		.out(chanx_right_out[10]));

	mux_2level_tapbuf_size3 mux_right_track_22 (
		.in({chany_top_in[13], chany_top_in[43], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_}),
		.sram(mux_2level_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_10_sram_inv[0:1]),
		.out(chanx_right_out[11]));

	mux_2level_tapbuf_size3 mux_right_track_24 (
		.in({chany_top_in[14], chany_top_in[47], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_11_sram_inv[0:1]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size3 mux_right_track_26 (
		.in({chany_top_in[16], chany_top_in[51], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_}),
		.sram(mux_2level_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_12_sram_inv[0:1]),
		.out(chanx_right_out[13]));

	mux_2level_tapbuf_size3 mux_right_track_28 (
		.in({chany_top_in[17], chany_top_in[55], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_}),
		.sram(mux_2level_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_13_sram_inv[0:1]),
		.out(chanx_right_out[14]));

	mux_2level_tapbuf_size3 mux_right_track_30 (
		.in({chany_top_in[18], chany_top_in[59], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_}),
		.sram(mux_2level_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_14_sram_inv[0:1]),
		.out(chanx_right_out[15]));

	mux_2level_tapbuf_size3 mux_right_track_32 (
		.in({chany_top_in[20], chany_top_in[63], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_15_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size3 mux_right_track_34 (
		.in({chany_top_in[21], chany_top_in[67], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_}),
		.sram(mux_2level_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_16_sram_inv[0:1]),
		.out(chanx_right_out[17]));

	mux_2level_tapbuf_size3 mux_right_track_36 (
		.in({chany_top_in[22], chany_top_in[71], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_17_sram_inv[0:1]),
		.out(chanx_right_out[18]));

	mux_2level_tapbuf_size3 mux_right_track_38 (
		.in({chany_top_in[24], chany_top_in[75], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_18_sram_inv[0:1]),
		.out(chanx_right_out[19]));

	mux_2level_tapbuf_size3 mux_right_track_40 (
		.in({chany_top_in[25], chany_top_in[79], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_}),
		.sram(mux_2level_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_19_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size3 mux_right_track_42 (
		.in({chany_top_in[26], chany_top_in[83], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_}),
		.sram(mux_2level_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_20_sram_inv[0:1]),
		.out(chanx_right_out[21]));

	mux_2level_tapbuf_size3 mux_right_track_44 (
		.in({chany_top_in[28], chany_top_in[87], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_21_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_2level_tapbuf_size3 mux_right_track_46 (
		.in({chany_top_in[29], chany_top_in[91], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_}),
		.sram(mux_2level_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_22_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_2level_tapbuf_size3 mux_right_track_48 (
		.in({chany_top_in[30], chany_top_in[95], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_}),
		.sram(mux_2level_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_23_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size3 mux_right_track_50 (
		.in({chany_top_in[32], chany_top_in[99], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_}),
		.sram(mux_2level_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_24_sram_inv[0:1]),
		.out(chanx_right_out[25]));

	mux_2level_tapbuf_size3 mux_right_track_52 (
		.in({chany_top_in[33], chany_top_in[103], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_25_sram_inv[0:1]),
		.out(chanx_right_out[26]));

	mux_2level_tapbuf_size3 mux_right_track_54 (
		.in({chany_top_in[34], chany_top_in[107], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_}),
		.sram(mux_2level_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_26_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_2level_tapbuf_size3 mux_right_track_56 (
		.in({chany_top_in[36], chany_top_in[111], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_27_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_2level_tapbuf_size3 mux_right_track_58 (
		.in({chany_top_in[37], chany_top_in[115], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_28_sram_inv[0:1]),
		.out(chanx_right_out[29]));

	mux_2level_tapbuf_size3 mux_right_track_60 (
		.in({chany_top_in[38], chany_top_in[119], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_}),
		.sram(mux_2level_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_29_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_2level_tapbuf_size3 mux_right_track_62 (
		.in({chany_top_in[40], chany_top_in[123], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_}),
		.sram(mux_2level_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_30_sram_inv[0:1]),
		.out(chanx_right_out[31]));

	mux_2level_tapbuf_size3 mux_right_track_64 (
		.in({chany_top_in[41], chany_top_in[127], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_31_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size3 mux_right_track_66 (
		.in({chany_top_in[42], chany_top_in[131], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_}),
		.sram(mux_2level_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_32_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	mux_2level_tapbuf_size3 mux_right_track_68 (
		.in({chany_top_in[44], chany_top_in[135], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_}),
		.sram(mux_2level_tapbuf_size3_33_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_33_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_2level_tapbuf_size3 mux_right_track_70 (
		.in({chany_top_in[45], chany_top_in[139], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_}),
		.sram(mux_2level_tapbuf_size3_34_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_34_sram_inv[0:1]),
		.out(chanx_right_out[35]));

	mux_2level_tapbuf_size3 mux_right_track_72 (
		.in({chany_top_in[46], chany_top_in[143], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size3_35_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_35_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size3 mux_right_track_78 (
		.in({chany_top_in[50], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chany_bottom_in[145]}),
		.sram(mux_2level_tapbuf_size3_36_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_36_sram_inv[0:1]),
		.out(chanx_right_out[39]));

	mux_2level_tapbuf_size3 mux_right_track_80 (
		.in({chany_top_in[52], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[144]}),
		.sram(mux_2level_tapbuf_size3_37_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_37_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size3 mux_right_track_82 (
		.in({chany_top_in[53], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[142]}),
		.sram(mux_2level_tapbuf_size3_38_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_38_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	mux_2level_tapbuf_size3 mux_right_track_84 (
		.in({chany_top_in[54], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[141]}),
		.sram(mux_2level_tapbuf_size3_39_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_39_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_2level_tapbuf_size3 mux_right_track_86 (
		.in({chany_top_in[56], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, chany_bottom_in[140]}),
		.sram(mux_2level_tapbuf_size3_40_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_40_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_2level_tapbuf_size3 mux_right_track_88 (
		.in({chany_top_in[57], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[138]}),
		.sram(mux_2level_tapbuf_size3_41_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_41_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	mux_2level_tapbuf_size3 mux_right_track_90 (
		.in({chany_top_in[58], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[137]}),
		.sram(mux_2level_tapbuf_size3_42_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_42_sram_inv[0:1]),
		.out(chanx_right_out[45]));

	mux_2level_tapbuf_size3 mux_right_track_92 (
		.in({chany_top_in[60], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[136]}),
		.sram(mux_2level_tapbuf_size3_43_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_43_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	mux_2level_tapbuf_size3 mux_right_track_94 (
		.in({chany_top_in[61], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[134]}),
		.sram(mux_2level_tapbuf_size3_44_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_44_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_2level_tapbuf_size3 mux_right_track_96 (
		.in({chany_top_in[62], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[133]}),
		.sram(mux_2level_tapbuf_size3_45_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_45_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_2level_tapbuf_size3 mux_right_track_98 (
		.in({chany_top_in[64], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chany_bottom_in[132]}),
		.sram(mux_2level_tapbuf_size3_46_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_46_sram_inv[0:1]),
		.out(chanx_right_out[49]));

	mux_2level_tapbuf_size3 mux_right_track_100 (
		.in({chany_top_in[65], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[130]}),
		.sram(mux_2level_tapbuf_size3_47_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_47_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	mux_2level_tapbuf_size3 mux_right_track_102 (
		.in({chany_top_in[66], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[129]}),
		.sram(mux_2level_tapbuf_size3_48_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_48_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	mux_2level_tapbuf_size3 mux_right_track_104 (
		.in({chany_top_in[68], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[128]}),
		.sram(mux_2level_tapbuf_size3_49_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_49_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	mux_2level_tapbuf_size3 mux_right_track_106 (
		.in({chany_top_in[69], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, chany_bottom_in[126]}),
		.sram(mux_2level_tapbuf_size3_50_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_50_sram_inv[0:1]),
		.out(chanx_right_out[53]));

	mux_2level_tapbuf_size3 mux_right_track_108 (
		.in({chany_top_in[70], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[125]}),
		.sram(mux_2level_tapbuf_size3_51_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_51_sram_inv[0:1]),
		.out(chanx_right_out[54]));

	mux_2level_tapbuf_size3 mux_right_track_110 (
		.in({chany_top_in[72], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[124]}),
		.sram(mux_2level_tapbuf_size3_52_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_52_sram_inv[0:1]),
		.out(chanx_right_out[55]));

	mux_2level_tapbuf_size3 mux_right_track_112 (
		.in({chany_top_in[73], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[122]}),
		.sram(mux_2level_tapbuf_size3_53_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_53_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_2level_tapbuf_size3 mux_right_track_114 (
		.in({chany_top_in[74], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[121]}),
		.sram(mux_2level_tapbuf_size3_54_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_54_sram_inv[0:1]),
		.out(chanx_right_out[57]));

	mux_2level_tapbuf_size3 mux_right_track_116 (
		.in({chany_top_in[76], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[120]}),
		.sram(mux_2level_tapbuf_size3_55_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_55_sram_inv[0:1]),
		.out(chanx_right_out[58]));

	mux_2level_tapbuf_size3 mux_right_track_118 (
		.in({chany_top_in[77], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chany_bottom_in[118]}),
		.sram(mux_2level_tapbuf_size3_56_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_56_sram_inv[0:1]),
		.out(chanx_right_out[59]));

	mux_2level_tapbuf_size3 mux_right_track_120 (
		.in({chany_top_in[78], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[117]}),
		.sram(mux_2level_tapbuf_size3_57_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_57_sram_inv[0:1]),
		.out(chanx_right_out[60]));

	mux_2level_tapbuf_size3 mux_right_track_122 (
		.in({chany_top_in[80], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[116]}),
		.sram(mux_2level_tapbuf_size3_58_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_58_sram_inv[0:1]),
		.out(chanx_right_out[61]));

	mux_2level_tapbuf_size3 mux_right_track_124 (
		.in({chany_top_in[81], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[114]}),
		.sram(mux_2level_tapbuf_size3_59_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_59_sram_inv[0:1]),
		.out(chanx_right_out[62]));

	mux_2level_tapbuf_size3 mux_right_track_126 (
		.in({chany_top_in[82], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, chany_bottom_in[113]}),
		.sram(mux_2level_tapbuf_size3_60_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_60_sram_inv[0:1]),
		.out(chanx_right_out[63]));

	mux_2level_tapbuf_size3 mux_right_track_128 (
		.in({chany_top_in[84], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[112]}),
		.sram(mux_2level_tapbuf_size3_61_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_61_sram_inv[0:1]),
		.out(chanx_right_out[64]));

	mux_2level_tapbuf_size3 mux_right_track_130 (
		.in({chany_top_in[85], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[110]}),
		.sram(mux_2level_tapbuf_size3_62_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_62_sram_inv[0:1]),
		.out(chanx_right_out[65]));

	mux_2level_tapbuf_size3 mux_right_track_132 (
		.in({chany_top_in[86], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[109]}),
		.sram(mux_2level_tapbuf_size3_63_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_63_sram_inv[0:1]),
		.out(chanx_right_out[66]));

	mux_2level_tapbuf_size3 mux_right_track_134 (
		.in({chany_top_in[88], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[108]}),
		.sram(mux_2level_tapbuf_size3_64_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_64_sram_inv[0:1]),
		.out(chanx_right_out[67]));

	mux_2level_tapbuf_size3 mux_right_track_136 (
		.in({chany_top_in[89], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[106]}),
		.sram(mux_2level_tapbuf_size3_65_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_65_sram_inv[0:1]),
		.out(chanx_right_out[68]));

	mux_2level_tapbuf_size3 mux_right_track_138 (
		.in({chany_top_in[90], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chany_bottom_in[105]}),
		.sram(mux_2level_tapbuf_size3_66_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_66_sram_inv[0:1]),
		.out(chanx_right_out[69]));

	mux_2level_tapbuf_size3 mux_right_track_140 (
		.in({chany_top_in[92], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[104]}),
		.sram(mux_2level_tapbuf_size3_67_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_67_sram_inv[0:1]),
		.out(chanx_right_out[70]));

	mux_2level_tapbuf_size3 mux_right_track_142 (
		.in({chany_top_in[93], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[102]}),
		.sram(mux_2level_tapbuf_size3_68_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_68_sram_inv[0:1]),
		.out(chanx_right_out[71]));

	mux_2level_tapbuf_size3 mux_right_track_144 (
		.in({chany_top_in[94], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[101]}),
		.sram(mux_2level_tapbuf_size3_69_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_69_sram_inv[0:1]),
		.out(chanx_right_out[72]));

	mux_2level_tapbuf_size3 mux_right_track_146 (
		.in({chany_top_in[96], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, chany_bottom_in[100]}),
		.sram(mux_2level_tapbuf_size3_70_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_70_sram_inv[0:1]),
		.out(chanx_right_out[73]));

	mux_2level_tapbuf_size3 mux_right_track_148 (
		.in({chany_top_in[97], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[98]}),
		.sram(mux_2level_tapbuf_size3_71_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_71_sram_inv[0:1]),
		.out(chanx_right_out[74]));

	mux_2level_tapbuf_size3 mux_right_track_150 (
		.in({chany_top_in[98], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[97]}),
		.sram(mux_2level_tapbuf_size3_72_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_72_sram_inv[0:1]),
		.out(chanx_right_out[75]));

	mux_2level_tapbuf_size3 mux_right_track_152 (
		.in({chany_top_in[100], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[96]}),
		.sram(mux_2level_tapbuf_size3_73_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_73_sram_inv[0:1]),
		.out(chanx_right_out[76]));

	mux_2level_tapbuf_size3 mux_right_track_154 (
		.in({chany_top_in[101], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[94]}),
		.sram(mux_2level_tapbuf_size3_74_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_74_sram_inv[0:1]),
		.out(chanx_right_out[77]));

	mux_2level_tapbuf_size3 mux_right_track_156 (
		.in({chany_top_in[102], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[93]}),
		.sram(mux_2level_tapbuf_size3_75_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_75_sram_inv[0:1]),
		.out(chanx_right_out[78]));

	mux_2level_tapbuf_size3 mux_right_track_158 (
		.in({chany_top_in[104], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chany_bottom_in[92]}),
		.sram(mux_2level_tapbuf_size3_76_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_76_sram_inv[0:1]),
		.out(chanx_right_out[79]));

	mux_2level_tapbuf_size3 mux_right_track_160 (
		.in({chany_top_in[105], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[90]}),
		.sram(mux_2level_tapbuf_size3_77_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_77_sram_inv[0:1]),
		.out(chanx_right_out[80]));

	mux_2level_tapbuf_size3 mux_right_track_162 (
		.in({chany_top_in[106], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[89]}),
		.sram(mux_2level_tapbuf_size3_78_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_78_sram_inv[0:1]),
		.out(chanx_right_out[81]));

	mux_2level_tapbuf_size3 mux_right_track_164 (
		.in({chany_top_in[108], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[88]}),
		.sram(mux_2level_tapbuf_size3_79_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_79_sram_inv[0:1]),
		.out(chanx_right_out[82]));

	mux_2level_tapbuf_size3 mux_right_track_166 (
		.in({chany_top_in[109], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, chany_bottom_in[86]}),
		.sram(mux_2level_tapbuf_size3_80_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_80_sram_inv[0:1]),
		.out(chanx_right_out[83]));

	mux_2level_tapbuf_size3 mux_right_track_168 (
		.in({chany_top_in[110], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[85]}),
		.sram(mux_2level_tapbuf_size3_81_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_81_sram_inv[0:1]),
		.out(chanx_right_out[84]));

	mux_2level_tapbuf_size3 mux_right_track_170 (
		.in({chany_top_in[112], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[84]}),
		.sram(mux_2level_tapbuf_size3_82_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_82_sram_inv[0:1]),
		.out(chanx_right_out[85]));

	mux_2level_tapbuf_size3 mux_right_track_172 (
		.in({chany_top_in[113], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[82]}),
		.sram(mux_2level_tapbuf_size3_83_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_83_sram_inv[0:1]),
		.out(chanx_right_out[86]));

	mux_2level_tapbuf_size3 mux_right_track_174 (
		.in({chany_top_in[114], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[81]}),
		.sram(mux_2level_tapbuf_size3_84_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_84_sram_inv[0:1]),
		.out(chanx_right_out[87]));

	mux_2level_tapbuf_size3 mux_right_track_176 (
		.in({chany_top_in[116], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[80]}),
		.sram(mux_2level_tapbuf_size3_85_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_85_sram_inv[0:1]),
		.out(chanx_right_out[88]));

	mux_2level_tapbuf_size3 mux_right_track_178 (
		.in({chany_top_in[117], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chany_bottom_in[78]}),
		.sram(mux_2level_tapbuf_size3_86_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_86_sram_inv[0:1]),
		.out(chanx_right_out[89]));

	mux_2level_tapbuf_size3 mux_right_track_180 (
		.in({chany_top_in[118], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[77]}),
		.sram(mux_2level_tapbuf_size3_87_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_87_sram_inv[0:1]),
		.out(chanx_right_out[90]));

	mux_2level_tapbuf_size3 mux_right_track_182 (
		.in({chany_top_in[120], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[76]}),
		.sram(mux_2level_tapbuf_size3_88_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_88_sram_inv[0:1]),
		.out(chanx_right_out[91]));

	mux_2level_tapbuf_size3 mux_right_track_184 (
		.in({chany_top_in[121], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[74]}),
		.sram(mux_2level_tapbuf_size3_89_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_89_sram_inv[0:1]),
		.out(chanx_right_out[92]));

	mux_2level_tapbuf_size3 mux_right_track_186 (
		.in({chany_top_in[122], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, chany_bottom_in[73]}),
		.sram(mux_2level_tapbuf_size3_90_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_90_sram_inv[0:1]),
		.out(chanx_right_out[93]));

	mux_2level_tapbuf_size3 mux_right_track_188 (
		.in({chany_top_in[124], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[72]}),
		.sram(mux_2level_tapbuf_size3_91_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_91_sram_inv[0:1]),
		.out(chanx_right_out[94]));

	mux_2level_tapbuf_size3 mux_right_track_190 (
		.in({chany_top_in[125], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[70]}),
		.sram(mux_2level_tapbuf_size3_92_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_92_sram_inv[0:1]),
		.out(chanx_right_out[95]));

	mux_2level_tapbuf_size3 mux_right_track_192 (
		.in({chany_top_in[126], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[69]}),
		.sram(mux_2level_tapbuf_size3_93_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_93_sram_inv[0:1]),
		.out(chanx_right_out[96]));

	mux_2level_tapbuf_size3 mux_right_track_194 (
		.in({chany_top_in[128], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[68]}),
		.sram(mux_2level_tapbuf_size3_94_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_94_sram_inv[0:1]),
		.out(chanx_right_out[97]));

	mux_2level_tapbuf_size3 mux_right_track_196 (
		.in({chany_top_in[129], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[66]}),
		.sram(mux_2level_tapbuf_size3_95_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_95_sram_inv[0:1]),
		.out(chanx_right_out[98]));

	mux_2level_tapbuf_size3 mux_right_track_198 (
		.in({chany_top_in[130], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chany_bottom_in[65]}),
		.sram(mux_2level_tapbuf_size3_96_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_96_sram_inv[0:1]),
		.out(chanx_right_out[99]));

	mux_2level_tapbuf_size3 mux_right_track_200 (
		.in({chany_top_in[132], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[64]}),
		.sram(mux_2level_tapbuf_size3_97_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_97_sram_inv[0:1]),
		.out(chanx_right_out[100]));

	mux_2level_tapbuf_size3 mux_right_track_202 (
		.in({chany_top_in[133], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[62]}),
		.sram(mux_2level_tapbuf_size3_98_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_98_sram_inv[0:1]),
		.out(chanx_right_out[101]));

	mux_2level_tapbuf_size3 mux_right_track_204 (
		.in({chany_top_in[134], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[61]}),
		.sram(mux_2level_tapbuf_size3_99_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_99_sram_inv[0:1]),
		.out(chanx_right_out[102]));

	mux_2level_tapbuf_size3 mux_right_track_206 (
		.in({chany_top_in[136], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, chany_bottom_in[60]}),
		.sram(mux_2level_tapbuf_size3_100_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_100_sram_inv[0:1]),
		.out(chanx_right_out[103]));

	mux_2level_tapbuf_size3 mux_right_track_208 (
		.in({chany_top_in[137], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[58]}),
		.sram(mux_2level_tapbuf_size3_101_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_101_sram_inv[0:1]),
		.out(chanx_right_out[104]));

	mux_2level_tapbuf_size3 mux_right_track_210 (
		.in({chany_top_in[138], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[57]}),
		.sram(mux_2level_tapbuf_size3_102_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_102_sram_inv[0:1]),
		.out(chanx_right_out[105]));

	mux_2level_tapbuf_size3 mux_right_track_212 (
		.in({chany_top_in[140], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[56]}),
		.sram(mux_2level_tapbuf_size3_103_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_103_sram_inv[0:1]),
		.out(chanx_right_out[106]));

	mux_2level_tapbuf_size3 mux_right_track_214 (
		.in({chany_top_in[141], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[54]}),
		.sram(mux_2level_tapbuf_size3_104_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_104_sram_inv[0:1]),
		.out(chanx_right_out[107]));

	mux_2level_tapbuf_size3 mux_right_track_216 (
		.in({chany_top_in[142], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[53]}),
		.sram(mux_2level_tapbuf_size3_105_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_105_sram_inv[0:1]),
		.out(chanx_right_out[108]));

	mux_2level_tapbuf_size3 mux_right_track_218 (
		.in({chany_top_in[144], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chany_bottom_in[52]}),
		.sram(mux_2level_tapbuf_size3_106_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_106_sram_inv[0:1]),
		.out(chanx_right_out[109]));

	mux_2level_tapbuf_size3 mux_right_track_220 (
		.in({chany_top_in[145], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[50]}),
		.sram(mux_2level_tapbuf_size3_107_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_107_sram_inv[0:1]),
		.out(chanx_right_out[110]));

	mux_2level_tapbuf_size3 mux_right_track_226 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, chany_bottom_in[46], chany_bottom_in[143]}),
		.sram(mux_2level_tapbuf_size3_108_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_108_sram_inv[0:1]),
		.out(chanx_right_out[113]));

	mux_2level_tapbuf_size3 mux_right_track_228 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[45], chany_bottom_in[139]}),
		.sram(mux_2level_tapbuf_size3_109_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_109_sram_inv[0:1]),
		.out(chanx_right_out[114]));

	mux_2level_tapbuf_size3 mux_right_track_230 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[44], chany_bottom_in[135]}),
		.sram(mux_2level_tapbuf_size3_110_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_110_sram_inv[0:1]),
		.out(chanx_right_out[115]));

	mux_2level_tapbuf_size3 mux_right_track_232 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[42], chany_bottom_in[131]}),
		.sram(mux_2level_tapbuf_size3_111_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_111_sram_inv[0:1]),
		.out(chanx_right_out[116]));

	mux_2level_tapbuf_size3 mux_right_track_234 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[41], chany_bottom_in[127]}),
		.sram(mux_2level_tapbuf_size3_112_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_112_sram_inv[0:1]),
		.out(chanx_right_out[117]));

	mux_2level_tapbuf_size3 mux_right_track_236 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[40], chany_bottom_in[123]}),
		.sram(mux_2level_tapbuf_size3_113_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_113_sram_inv[0:1]),
		.out(chanx_right_out[118]));

	mux_2level_tapbuf_size3 mux_right_track_238 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chany_bottom_in[38], chany_bottom_in[119]}),
		.sram(mux_2level_tapbuf_size3_114_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_114_sram_inv[0:1]),
		.out(chanx_right_out[119]));

	mux_2level_tapbuf_size3 mux_right_track_240 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[37], chany_bottom_in[115]}),
		.sram(mux_2level_tapbuf_size3_115_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_115_sram_inv[0:1]),
		.out(chanx_right_out[120]));

	mux_2level_tapbuf_size3 mux_right_track_242 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[36], chany_bottom_in[111]}),
		.sram(mux_2level_tapbuf_size3_116_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_116_sram_inv[0:1]),
		.out(chanx_right_out[121]));

	mux_2level_tapbuf_size3 mux_right_track_244 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[34], chany_bottom_in[107]}),
		.sram(mux_2level_tapbuf_size3_117_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_117_sram_inv[0:1]),
		.out(chanx_right_out[122]));

	mux_2level_tapbuf_size3 mux_right_track_246 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, chany_bottom_in[33], chany_bottom_in[103]}),
		.sram(mux_2level_tapbuf_size3_118_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_118_sram_inv[0:1]),
		.out(chanx_right_out[123]));

	mux_2level_tapbuf_size3 mux_right_track_248 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[32], chany_bottom_in[99]}),
		.sram(mux_2level_tapbuf_size3_119_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_119_sram_inv[0:1]),
		.out(chanx_right_out[124]));

	mux_2level_tapbuf_size3 mux_right_track_250 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[30], chany_bottom_in[95]}),
		.sram(mux_2level_tapbuf_size3_120_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_120_sram_inv[0:1]),
		.out(chanx_right_out[125]));

	mux_2level_tapbuf_size3 mux_right_track_252 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[29], chany_bottom_in[91]}),
		.sram(mux_2level_tapbuf_size3_121_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_121_sram_inv[0:1]),
		.out(chanx_right_out[126]));

	mux_2level_tapbuf_size3 mux_right_track_254 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[28], chany_bottom_in[87]}),
		.sram(mux_2level_tapbuf_size3_122_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_122_sram_inv[0:1]),
		.out(chanx_right_out[127]));

	mux_2level_tapbuf_size3 mux_right_track_256 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[26], chany_bottom_in[83]}),
		.sram(mux_2level_tapbuf_size3_123_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_123_sram_inv[0:1]),
		.out(chanx_right_out[128]));

	mux_2level_tapbuf_size3 mux_right_track_258 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chany_bottom_in[25], chany_bottom_in[79]}),
		.sram(mux_2level_tapbuf_size3_124_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_124_sram_inv[0:1]),
		.out(chanx_right_out[129]));

	mux_2level_tapbuf_size3 mux_right_track_260 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[24], chany_bottom_in[75]}),
		.sram(mux_2level_tapbuf_size3_125_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_125_sram_inv[0:1]),
		.out(chanx_right_out[130]));

	mux_2level_tapbuf_size3 mux_right_track_262 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[22], chany_bottom_in[71]}),
		.sram(mux_2level_tapbuf_size3_126_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_126_sram_inv[0:1]),
		.out(chanx_right_out[131]));

	mux_2level_tapbuf_size3 mux_right_track_264 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[21], chany_bottom_in[67]}),
		.sram(mux_2level_tapbuf_size3_127_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_127_sram_inv[0:1]),
		.out(chanx_right_out[132]));

	mux_2level_tapbuf_size3 mux_right_track_266 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, chany_bottom_in[20], chany_bottom_in[63]}),
		.sram(mux_2level_tapbuf_size3_128_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_128_sram_inv[0:1]),
		.out(chanx_right_out[133]));

	mux_2level_tapbuf_size3 mux_right_track_268 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[18], chany_bottom_in[59]}),
		.sram(mux_2level_tapbuf_size3_129_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_129_sram_inv[0:1]),
		.out(chanx_right_out[134]));

	mux_2level_tapbuf_size3 mux_right_track_270 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[17], chany_bottom_in[55]}),
		.sram(mux_2level_tapbuf_size3_130_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_130_sram_inv[0:1]),
		.out(chanx_right_out[135]));

	mux_2level_tapbuf_size3 mux_right_track_272 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[16], chany_bottom_in[51]}),
		.sram(mux_2level_tapbuf_size3_131_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_131_sram_inv[0:1]),
		.out(chanx_right_out[136]));

	mux_2level_tapbuf_size3 mux_right_track_274 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[14], chany_bottom_in[47]}),
		.sram(mux_2level_tapbuf_size3_132_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_132_sram_inv[0:1]),
		.out(chanx_right_out[137]));

	mux_2level_tapbuf_size3 mux_right_track_276 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[13], chany_bottom_in[43]}),
		.sram(mux_2level_tapbuf_size3_133_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_133_sram_inv[0:1]),
		.out(chanx_right_out[138]));

	mux_2level_tapbuf_size3 mux_right_track_278 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chany_bottom_in[12], chany_bottom_in[39]}),
		.sram(mux_2level_tapbuf_size3_134_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_134_sram_inv[0:1]),
		.out(chanx_right_out[139]));

	mux_2level_tapbuf_size3 mux_right_track_280 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[10], chany_bottom_in[35]}),
		.sram(mux_2level_tapbuf_size3_135_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_135_sram_inv[0:1]),
		.out(chanx_right_out[140]));

	mux_2level_tapbuf_size3 mux_right_track_282 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[9], chany_bottom_in[31]}),
		.sram(mux_2level_tapbuf_size3_136_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_136_sram_inv[0:1]),
		.out(chanx_right_out[141]));

	mux_2level_tapbuf_size3 mux_right_track_284 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[8], chany_bottom_in[27]}),
		.sram(mux_2level_tapbuf_size3_137_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_137_sram_inv[0:1]),
		.out(chanx_right_out[142]));

	mux_2level_tapbuf_size3 mux_right_track_286 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, chany_bottom_in[6], chany_bottom_in[23]}),
		.sram(mux_2level_tapbuf_size3_138_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_138_sram_inv[0:1]),
		.out(chanx_right_out[143]));

	mux_2level_tapbuf_size3 mux_right_track_288 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[5], chany_bottom_in[19]}),
		.sram(mux_2level_tapbuf_size3_139_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_139_sram_inv[0:1]),
		.out(chanx_right_out[144]));

	mux_2level_tapbuf_size3 mux_right_track_290 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[4], chany_bottom_in[15]}),
		.sram(mux_2level_tapbuf_size3_140_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_140_sram_inv[0:1]),
		.out(chanx_right_out[145]));

	mux_2level_tapbuf_size3 mux_right_track_292 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[2], chany_bottom_in[11]}),
		.sram(mux_2level_tapbuf_size3_141_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_141_sram_inv[0:1]),
		.out(chanx_right_out[146]));

	mux_2level_tapbuf_size3 mux_right_track_294 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[1], chany_bottom_in[7]}),
		.sram(mux_2level_tapbuf_size3_142_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_142_sram_inv[0:1]),
		.out(chanx_right_out[147]));

	mux_2level_tapbuf_size3 mux_right_track_296 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[0], chany_bottom_in[3]}),
		.sram(mux_2level_tapbuf_size3_143_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_143_sram_inv[0:1]),
		.out(chanx_right_out[148]));

	mux_2level_tapbuf_size3_mem mem_right_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_0_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_1_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_6 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_2_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_3_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_4_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_5_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_14 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_6_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_7_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_8_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_9_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_22 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_10_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_11_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_12_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_13_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_30 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_14_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_15_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_34 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_16_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_17_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_38 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_18_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_19_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_20_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_21_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_46 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_22_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_23_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_24_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_52 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_25_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_54 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_26_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_27_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_28_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_29_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_62 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_30_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_31_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_32_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_33_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_33_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_70 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_34_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_34_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_35_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_35_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_78 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_36_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_36_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_37_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_37_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_38_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_38_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_39_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_39_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_86 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_40_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_40_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_41_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_41_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_42_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_42_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_43_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_43_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_94 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_44_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_44_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_45_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_45_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_46_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_46_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_47_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_47_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_102 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_48_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_48_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_49_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_49_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_106 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_50_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_50_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_51_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_51_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_110 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_52_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_52_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_53_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_53_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_54_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_54_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_55_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_55_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_118 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_56_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_56_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_57_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_57_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_58_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_58_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_124 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_59_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_59_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_126 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_60_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_60_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_61_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_61_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_62_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_62_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_63_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_63_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_134 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_64_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_64_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_65_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_65_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_138 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_66_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_66_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_67_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_67_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_142 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_68_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_68_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_69_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_69_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_70_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_70_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_71_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_71_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_150 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_72_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_72_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_73_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_73_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_74_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_74_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_75_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_75_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_158 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_76_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_76_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_77_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_77_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_78_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_78_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_78_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_79_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_79_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_79_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_166 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_79_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_80_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_80_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_80_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_80_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_81_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_81_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_81_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_81_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_82_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_82_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_82_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_82_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_83_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_83_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_83_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_174 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_83_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_84_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_84_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_84_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_84_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_85_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_85_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_85_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_178 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_85_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_86_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_86_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_86_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_86_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_87_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_87_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_87_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_182 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_87_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_88_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_88_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_88_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_88_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_89_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_89_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_89_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_89_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_90_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_90_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_90_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_90_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_91_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_91_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_91_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_190 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_91_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_92_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_92_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_92_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_92_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_93_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_93_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_93_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_93_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_94_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_94_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_94_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_196 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_94_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_95_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_95_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_95_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_198 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_95_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_96_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_96_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_96_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_96_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_97_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_97_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_97_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_97_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_98_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_98_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_98_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_98_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_99_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_99_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_99_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_206 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_99_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_100_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_100_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_100_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_100_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_101_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_101_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_101_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_210 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_101_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_102_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_102_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_102_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_212 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_102_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_103_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_103_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_103_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_214 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_103_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_104_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_104_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_104_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_104_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_105_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_105_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_105_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_218 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_105_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_106_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_106_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_106_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_220 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_106_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_107_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_107_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_107_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_226 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_108_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_108_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_108_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_228 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_108_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_109_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_109_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_109_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_230 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_109_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_110_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_110_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_110_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_110_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_111_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_111_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_111_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_234 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_111_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_112_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_112_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_112_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_236 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_112_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_113_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_113_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_113_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_238 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_113_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_114_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_114_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_114_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_114_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_115_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_115_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_115_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_242 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_115_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_116_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_116_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_116_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_244 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_116_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_117_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_117_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_117_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_246 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_117_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_118_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_118_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_118_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_118_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_119_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_119_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_119_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_250 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_119_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_120_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_120_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_120_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_252 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_120_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_121_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_121_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_121_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_254 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_121_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_122_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_122_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_122_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_122_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_123_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_123_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_123_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_258 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_123_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_124_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_124_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_124_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_260 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_124_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_125_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_125_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_125_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_262 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_125_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_126_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_126_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_126_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_126_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_127_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_127_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_127_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_266 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_127_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_128_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_128_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_128_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_268 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_128_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_129_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_129_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_129_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_270 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_129_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_130_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_130_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_130_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_130_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_131_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_131_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_131_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_274 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_131_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_132_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_132_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_132_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_276 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_132_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_133_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_133_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_133_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_278 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_133_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_134_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_134_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_134_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_134_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_135_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_135_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_135_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_282 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_135_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_136_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_136_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_136_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_284 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_136_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_137_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_137_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_137_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_286 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_137_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_138_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_138_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_138_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_138_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_139_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_139_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_139_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_290 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_139_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_140_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_140_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_140_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_292 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_140_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_141_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_141_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_141_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_294 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_141_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_142_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_142_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_142_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_142_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_143_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_143_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_143_sram_inv[0:1]));

	mux_2level_tapbuf_size4 mux_right_track_74 (
		.in({chany_top_in[48], chany_top_in[147], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, chany_bottom_in[148]}),
		.sram(mux_2level_tapbuf_size4_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_0_sram_inv[0:5]),
		.out(chanx_right_out[37]));

	mux_2level_tapbuf_size4 mux_right_track_76 (
		.in({chany_top_in[49], chany_top_in[149], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[146]}),
		.sram(mux_2level_tapbuf_size4_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_1_sram_inv[0:5]),
		.out(chanx_right_out[38]));

	mux_2level_tapbuf_size4 mux_right_track_222 (
		.in({chany_top_in[146], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[49], chany_bottom_in[149]}),
		.sram(mux_2level_tapbuf_size4_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_2_sram_inv[0:5]),
		.out(chanx_right_out[111]));

	mux_2level_tapbuf_size4 mux_right_track_224 (
		.in({chany_top_in[148], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[48], chany_bottom_in[147]}),
		.sram(mux_2level_tapbuf_size4_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_3_sram_inv[0:5]),
		.out(chanx_right_out[112]));

	mux_2level_tapbuf_size4_mem mem_right_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_0_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_1_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_222 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_107_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_2_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_3_sram_inv[0:5]));

	mux_2level_tapbuf_size11 mux_bottom_track_1 (
		.in({chany_top_in[0], chany_top_in[50], chany_top_in[101], chanx_right_in[36], chanx_right_in[74], chanx_right_in[112], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_29_}),
		.sram(mux_2level_tapbuf_size11_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_0_sram_inv[0:7]),
		.out(chany_bottom_out[0]));

	mux_2level_tapbuf_size11 mux_bottom_track_57 (
		.in({chany_top_in[9], chany_top_in[60], chany_top_in[110], chanx_right_in[29], chanx_right_in[67], chanx_right_in[105], chanx_right_in[143], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_27_}),
		.sram(mux_2level_tapbuf_size11_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_1_sram_inv[0:7]),
		.out(chany_bottom_out[28]));

	mux_2level_tapbuf_size11 mux_bottom_track_65 (
		.in({chany_top_in[10], chany_top_in[61], chany_top_in[112], chanx_right_in[28], chanx_right_in[66], chanx_right_in[104], chanx_right_in[142], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_28_}),
		.sram(mux_2level_tapbuf_size11_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_2_sram_inv[0:7]),
		.out(chany_bottom_out[32]));

	mux_2level_tapbuf_size11 mux_bottom_track_129 (
		.in({chany_top_in[21], chany_top_in[72], chany_top_in[122], chanx_right_in[20], chanx_right_in[58], chanx_right_in[96], chanx_right_in[134], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_27_}),
		.sram(mux_2level_tapbuf_size11_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_3_sram_inv[0:7]),
		.out(chany_bottom_out[64]));

	mux_2level_tapbuf_size11 mux_bottom_track_137 (
		.in({chany_top_in[22], chany_top_in[73], chany_top_in[124], chanx_right_in[19], chanx_right_in[57], chanx_right_in[95], chanx_right_in[133], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_28_}),
		.sram(mux_2level_tapbuf_size11_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_4_sram_inv[0:7]),
		.out(chany_bottom_out[68]));

	mux_2level_tapbuf_size11 mux_bottom_track_201 (
		.in({chany_top_in[33], chany_top_in[84], chany_top_in[134], chanx_right_in[11], chanx_right_in[49], chanx_right_in[87], chanx_right_in[125], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_27_}),
		.sram(mux_2level_tapbuf_size11_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_5_sram_inv[0:7]),
		.out(chany_bottom_out[100]));

	mux_2level_tapbuf_size11 mux_bottom_track_209 (
		.in({chany_top_in[34], chany_top_in[85], chany_top_in[136], chanx_right_in[10], chanx_right_in[48], chanx_right_in[86], chanx_right_in[124], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_28_}),
		.sram(mux_2level_tapbuf_size11_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_6_sram_inv[0:7]),
		.out(chany_bottom_out[104]));

	mux_2level_tapbuf_size11 mux_bottom_track_273 (
		.in({chany_top_in[45], chany_top_in[96], chany_top_in[146], chanx_right_in[2], chanx_right_in[40], chanx_right_in[78], chanx_right_in[116], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_34_}),
		.sram(mux_2level_tapbuf_size11_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_7_sram_inv[0:7]),
		.out(chany_bottom_out[136]));

	mux_2level_tapbuf_size11 mux_bottom_track_281 (
		.in({chany_top_in[46], chany_top_in[97], chany_top_in[148], chanx_right_in[1], chanx_right_in[39], chanx_right_in[77], chanx_right_in[115], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_35_}),
		.sram(mux_2level_tapbuf_size11_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_8_sram_inv[0:7]),
		.out(chany_bottom_out[140]));

	mux_2level_tapbuf_size11_mem mem_bottom_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_143_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_0_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_bottom_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_1_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_bottom_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_2_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_bottom_track_129 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_3_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_bottom_track_137 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_4_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_bottom_track_201 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_5_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_bottom_track_209 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_6_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_bottom_track_273 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_7_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_bottom_track_281 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_8_sram_inv[0:7]));

	mux_2level_tapbuf_size12 mux_bottom_track_9 (
		.in({chany_top_in[1], chany_top_in[52], chany_top_in[102], chanx_right_in[35], chanx_right_in[73], chanx_right_in[111], chanx_right_in[149], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_30_}),
		.sram(mux_2level_tapbuf_size12_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_0_sram_inv[0:7]),
		.out(chany_bottom_out[4]));

	mux_2level_tapbuf_size12 mux_bottom_track_17 (
		.in({chany_top_in[2], chany_top_in[53], chany_top_in[104], chanx_right_in[34], chanx_right_in[72], chanx_right_in[110], chanx_right_in[148], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_31_}),
		.sram(mux_2level_tapbuf_size12_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_1_sram_inv[0:7]),
		.out(chany_bottom_out[8]));

	mux_2level_tapbuf_size12 mux_bottom_track_25 (
		.in({chany_top_in[4], chany_top_in[54], chany_top_in[105], chanx_right_in[33], chanx_right_in[71], chanx_right_in[109], chanx_right_in[147], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_32_}),
		.sram(mux_2level_tapbuf_size12_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_2_sram_inv[0:7]),
		.out(chany_bottom_out[12]));

	mux_2level_tapbuf_size12 mux_bottom_track_33 (
		.in({chany_top_in[5], chany_top_in[56], chany_top_in[106], chanx_right_in[32], chanx_right_in[70], chanx_right_in[108], chanx_right_in[146], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_33_}),
		.sram(mux_2level_tapbuf_size12_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_3_sram_inv[0:7]),
		.out(chany_bottom_out[16]));

	mux_2level_tapbuf_size12 mux_bottom_track_41 (
		.in({chany_top_in[6], chany_top_in[57], chany_top_in[108], chanx_right_in[31], chanx_right_in[69], chanx_right_in[107], chanx_right_in[145], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_34_}),
		.sram(mux_2level_tapbuf_size12_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_4_sram_inv[0:7]),
		.out(chany_bottom_out[20]));

	mux_2level_tapbuf_size12 mux_bottom_track_49 (
		.in({chany_top_in[8], chany_top_in[58], chany_top_in[109], chanx_right_in[30], chanx_right_in[68], chanx_right_in[106], chanx_right_in[144], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_35_}),
		.sram(mux_2level_tapbuf_size12_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_5_sram_inv[0:7]),
		.out(chany_bottom_out[24]));

	mux_2level_tapbuf_size12 mux_bottom_track_73 (
		.in({chany_top_in[12], chany_top_in[62], chany_top_in[113], chanx_right_in[27], chanx_right_in[65], chanx_right_in[103], chanx_right_in[141], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_29_}),
		.sram(mux_2level_tapbuf_size12_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_6_sram_inv[0:7]),
		.out(chany_bottom_out[36]));

	mux_2level_tapbuf_size12 mux_bottom_track_81 (
		.in({chany_top_in[13], chany_top_in[64], chany_top_in[114], chanx_right_in[26], chanx_right_in[64], chanx_right_in[102], chanx_right_in[140], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_30_}),
		.sram(mux_2level_tapbuf_size12_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_7_sram_inv[0:7]),
		.out(chany_bottom_out[40]));

	mux_2level_tapbuf_size12 mux_bottom_track_89 (
		.in({chany_top_in[14], chany_top_in[65], chany_top_in[116], chanx_right_in[25], chanx_right_in[63], chanx_right_in[101], chanx_right_in[139], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_31_}),
		.sram(mux_2level_tapbuf_size12_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_8_sram_inv[0:7]),
		.out(chany_bottom_out[44]));

	mux_2level_tapbuf_size12 mux_bottom_track_97 (
		.in({chany_top_in[16], chany_top_in[66], chany_top_in[117], chanx_right_in[24], chanx_right_in[62], chanx_right_in[100], chanx_right_in[138], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_32_}),
		.sram(mux_2level_tapbuf_size12_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_9_sram_inv[0:7]),
		.out(chany_bottom_out[48]));

	mux_2level_tapbuf_size12 mux_bottom_track_105 (
		.in({chany_top_in[17], chany_top_in[68], chany_top_in[118], chanx_right_in[23], chanx_right_in[61], chanx_right_in[99], chanx_right_in[137], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_33_}),
		.sram(mux_2level_tapbuf_size12_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_10_sram_inv[0:7]),
		.out(chany_bottom_out[52]));

	mux_2level_tapbuf_size12 mux_bottom_track_113 (
		.in({chany_top_in[18], chany_top_in[69], chany_top_in[120], chanx_right_in[22], chanx_right_in[60], chanx_right_in[98], chanx_right_in[136], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_34_}),
		.sram(mux_2level_tapbuf_size12_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_11_sram_inv[0:7]),
		.out(chany_bottom_out[56]));

	mux_2level_tapbuf_size12 mux_bottom_track_121 (
		.in({chany_top_in[20], chany_top_in[70], chany_top_in[121], chanx_right_in[21], chanx_right_in[59], chanx_right_in[97], chanx_right_in[135], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_35_}),
		.sram(mux_2level_tapbuf_size12_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_12_sram_inv[0:7]),
		.out(chany_bottom_out[60]));

	mux_2level_tapbuf_size12 mux_bottom_track_145 (
		.in({chany_top_in[24], chany_top_in[74], chany_top_in[125], chanx_right_in[18], chanx_right_in[56], chanx_right_in[94], chanx_right_in[132], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_29_}),
		.sram(mux_2level_tapbuf_size12_13_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_13_sram_inv[0:7]),
		.out(chany_bottom_out[72]));

	mux_2level_tapbuf_size12 mux_bottom_track_153 (
		.in({chany_top_in[25], chany_top_in[76], chany_top_in[126], chanx_right_in[17], chanx_right_in[55], chanx_right_in[93], chanx_right_in[131], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_30_}),
		.sram(mux_2level_tapbuf_size12_14_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_14_sram_inv[0:7]),
		.out(chany_bottom_out[76]));

	mux_2level_tapbuf_size12 mux_bottom_track_161 (
		.in({chany_top_in[26], chany_top_in[77], chany_top_in[128], chanx_right_in[16], chanx_right_in[54], chanx_right_in[92], chanx_right_in[130], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_31_}),
		.sram(mux_2level_tapbuf_size12_15_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_15_sram_inv[0:7]),
		.out(chany_bottom_out[80]));

	mux_2level_tapbuf_size12 mux_bottom_track_169 (
		.in({chany_top_in[28], chany_top_in[78], chany_top_in[129], chanx_right_in[15], chanx_right_in[53], chanx_right_in[91], chanx_right_in[129], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_32_}),
		.sram(mux_2level_tapbuf_size12_16_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_16_sram_inv[0:7]),
		.out(chany_bottom_out[84]));

	mux_2level_tapbuf_size12 mux_bottom_track_177 (
		.in({chany_top_in[29], chany_top_in[80], chany_top_in[130], chanx_right_in[14], chanx_right_in[52], chanx_right_in[90], chanx_right_in[128], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_33_}),
		.sram(mux_2level_tapbuf_size12_17_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_17_sram_inv[0:7]),
		.out(chany_bottom_out[88]));

	mux_2level_tapbuf_size12 mux_bottom_track_185 (
		.in({chany_top_in[30], chany_top_in[81], chany_top_in[132], chanx_right_in[13], chanx_right_in[51], chanx_right_in[89], chanx_right_in[127], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_34_}),
		.sram(mux_2level_tapbuf_size12_18_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_18_sram_inv[0:7]),
		.out(chany_bottom_out[92]));

	mux_2level_tapbuf_size12 mux_bottom_track_193 (
		.in({chany_top_in[32], chany_top_in[82], chany_top_in[133], chanx_right_in[12], chanx_right_in[50], chanx_right_in[88], chanx_right_in[126], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_35_}),
		.sram(mux_2level_tapbuf_size12_19_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_19_sram_inv[0:7]),
		.out(chany_bottom_out[96]));

	mux_2level_tapbuf_size12 mux_bottom_track_217 (
		.in({chany_top_in[36], chany_top_in[86], chany_top_in[137], chanx_right_in[9], chanx_right_in[47], chanx_right_in[85], chanx_right_in[123], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_29_}),
		.sram(mux_2level_tapbuf_size12_20_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_20_sram_inv[0:7]),
		.out(chany_bottom_out[108]));

	mux_2level_tapbuf_size12 mux_bottom_track_225 (
		.in({chany_top_in[37], chany_top_in[88], chany_top_in[138], chanx_right_in[8], chanx_right_in[46], chanx_right_in[84], chanx_right_in[122], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_30_}),
		.sram(mux_2level_tapbuf_size12_21_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_21_sram_inv[0:7]),
		.out(chany_bottom_out[112]));

	mux_2level_tapbuf_size12 mux_bottom_track_233 (
		.in({chany_top_in[38], chany_top_in[89], chany_top_in[140], chanx_right_in[7], chanx_right_in[45], chanx_right_in[83], chanx_right_in[121], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_31_}),
		.sram(mux_2level_tapbuf_size12_22_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_22_sram_inv[0:7]),
		.out(chany_bottom_out[116]));

	mux_2level_tapbuf_size12 mux_bottom_track_241 (
		.in({chany_top_in[40], chany_top_in[90], chany_top_in[141], chanx_right_in[6], chanx_right_in[44], chanx_right_in[82], chanx_right_in[120], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_32_}),
		.sram(mux_2level_tapbuf_size12_23_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_23_sram_inv[0:7]),
		.out(chany_bottom_out[120]));

	mux_2level_tapbuf_size12 mux_bottom_track_249 (
		.in({chany_top_in[41], chany_top_in[92], chany_top_in[142], chanx_right_in[5], chanx_right_in[43], chanx_right_in[81], chanx_right_in[119], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_33_}),
		.sram(mux_2level_tapbuf_size12_24_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_24_sram_inv[0:7]),
		.out(chany_bottom_out[124]));

	mux_2level_tapbuf_size12 mux_bottom_track_257 (
		.in({chany_top_in[42], chany_top_in[93], chany_top_in[144], chanx_right_in[4], chanx_right_in[42], chanx_right_in[80], chanx_right_in[118], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_34_}),
		.sram(mux_2level_tapbuf_size12_25_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_25_sram_inv[0:7]),
		.out(chany_bottom_out[128]));

	mux_2level_tapbuf_size12 mux_bottom_track_265 (
		.in({chany_top_in[44], chany_top_in[94], chany_top_in[145], chanx_right_in[3], chanx_right_in[41], chanx_right_in[79], chanx_right_in[117], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_35_}),
		.sram(mux_2level_tapbuf_size12_26_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_26_sram_inv[0:7]),
		.out(chany_bottom_out[132]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_0_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_1_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_2_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_3_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_4_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_5_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_6_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_7_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_8_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_97 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_9_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_105 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_10_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_113 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_11_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_121 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_12_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_145 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_13_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_13_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_153 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_14_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_14_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_161 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_15_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_15_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_169 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_16_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_16_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_177 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_17_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_17_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_185 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_18_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_18_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_193 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_19_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_19_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_217 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_20_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_20_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_225 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_21_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_21_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_233 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_22_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_22_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_241 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_23_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_23_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_249 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_24_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_24_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_257 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_25_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_25_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_265 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_26_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_26_sram_inv[0:7]));

	mux_2level_tapbuf_size10 mux_bottom_track_289 (
		.in({chany_top_in[48], chany_top_in[98], chanx_right_in[0], chanx_right_in[38], chanx_right_in[76], chanx_right_in[114], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_27_}),
		.sram(mux_2level_tapbuf_size10_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_0_sram_inv[0:7]),
		.out(chany_bottom_out[144]));

	mux_2level_tapbuf_size10_mem mem_bottom_track_289 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_0_sram_inv[0:7]));

	mux_2level_tapbuf_size9 mux_bottom_track_297 (
		.in({chany_top_in[49], chany_top_in[100], chanx_right_in[37], chanx_right_in[75], chanx_right_in[113], bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_28_}),
		.sram(mux_2level_tapbuf_size9_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_0_sram_inv[0:7]),
		.out(chany_bottom_out[148]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_297 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_0_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_0_sram_inv[0:7]));

endmodule
// ----- END Verilog module for sb_6__1_ -----

//----- Default net type -----
`default_nettype wire



