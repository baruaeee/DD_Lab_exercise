//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][11]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Mon Jul  7 22:55:50 2025
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_0__11_ -----
module sb_0__11_(pReset,
                 prog_clk,
                 chanx_right_in,
                 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_,
                 chany_bottom_in,
                 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                 ccff_head,
                 chanx_right_out,
                 chany_bottom_out,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:149] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:149] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:149] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:149] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_2level_tapbuf_size2_0_sram;
wire [0:1] mux_2level_tapbuf_size2_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_100_sram;
wire [0:1] mux_2level_tapbuf_size2_100_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_101_sram;
wire [0:1] mux_2level_tapbuf_size2_101_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_102_sram;
wire [0:1] mux_2level_tapbuf_size2_102_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_103_sram;
wire [0:1] mux_2level_tapbuf_size2_103_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_104_sram;
wire [0:1] mux_2level_tapbuf_size2_104_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_105_sram;
wire [0:1] mux_2level_tapbuf_size2_105_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_106_sram;
wire [0:1] mux_2level_tapbuf_size2_106_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_107_sram;
wire [0:1] mux_2level_tapbuf_size2_107_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_108_sram;
wire [0:1] mux_2level_tapbuf_size2_108_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_109_sram;
wire [0:1] mux_2level_tapbuf_size2_109_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_10_sram;
wire [0:1] mux_2level_tapbuf_size2_10_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_110_sram;
wire [0:1] mux_2level_tapbuf_size2_110_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_111_sram;
wire [0:1] mux_2level_tapbuf_size2_111_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_112_sram;
wire [0:1] mux_2level_tapbuf_size2_112_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_113_sram;
wire [0:1] mux_2level_tapbuf_size2_113_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_114_sram;
wire [0:1] mux_2level_tapbuf_size2_114_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_115_sram;
wire [0:1] mux_2level_tapbuf_size2_115_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_116_sram;
wire [0:1] mux_2level_tapbuf_size2_116_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_117_sram;
wire [0:1] mux_2level_tapbuf_size2_117_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_118_sram;
wire [0:1] mux_2level_tapbuf_size2_118_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_119_sram;
wire [0:1] mux_2level_tapbuf_size2_119_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_11_sram;
wire [0:1] mux_2level_tapbuf_size2_11_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_120_sram;
wire [0:1] mux_2level_tapbuf_size2_120_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_121_sram;
wire [0:1] mux_2level_tapbuf_size2_121_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_122_sram;
wire [0:1] mux_2level_tapbuf_size2_122_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_123_sram;
wire [0:1] mux_2level_tapbuf_size2_123_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_124_sram;
wire [0:1] mux_2level_tapbuf_size2_124_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_125_sram;
wire [0:1] mux_2level_tapbuf_size2_125_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_126_sram;
wire [0:1] mux_2level_tapbuf_size2_126_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_127_sram;
wire [0:1] mux_2level_tapbuf_size2_127_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_128_sram;
wire [0:1] mux_2level_tapbuf_size2_128_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_129_sram;
wire [0:1] mux_2level_tapbuf_size2_129_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_12_sram;
wire [0:1] mux_2level_tapbuf_size2_12_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_130_sram;
wire [0:1] mux_2level_tapbuf_size2_130_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_131_sram;
wire [0:1] mux_2level_tapbuf_size2_131_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_132_sram;
wire [0:1] mux_2level_tapbuf_size2_132_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_133_sram;
wire [0:1] mux_2level_tapbuf_size2_133_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_134_sram;
wire [0:1] mux_2level_tapbuf_size2_134_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_135_sram;
wire [0:1] mux_2level_tapbuf_size2_135_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_136_sram;
wire [0:1] mux_2level_tapbuf_size2_136_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_137_sram;
wire [0:1] mux_2level_tapbuf_size2_137_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_138_sram;
wire [0:1] mux_2level_tapbuf_size2_138_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_139_sram;
wire [0:1] mux_2level_tapbuf_size2_139_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_13_sram;
wire [0:1] mux_2level_tapbuf_size2_13_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_140_sram;
wire [0:1] mux_2level_tapbuf_size2_140_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_141_sram;
wire [0:1] mux_2level_tapbuf_size2_141_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_142_sram;
wire [0:1] mux_2level_tapbuf_size2_142_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_143_sram;
wire [0:1] mux_2level_tapbuf_size2_143_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_144_sram;
wire [0:1] mux_2level_tapbuf_size2_144_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_145_sram;
wire [0:1] mux_2level_tapbuf_size2_145_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_146_sram;
wire [0:1] mux_2level_tapbuf_size2_146_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_147_sram;
wire [0:1] mux_2level_tapbuf_size2_147_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_148_sram;
wire [0:1] mux_2level_tapbuf_size2_148_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_149_sram;
wire [0:1] mux_2level_tapbuf_size2_149_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_14_sram;
wire [0:1] mux_2level_tapbuf_size2_14_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_150_sram;
wire [0:1] mux_2level_tapbuf_size2_150_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_151_sram;
wire [0:1] mux_2level_tapbuf_size2_151_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_152_sram;
wire [0:1] mux_2level_tapbuf_size2_152_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_153_sram;
wire [0:1] mux_2level_tapbuf_size2_153_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_154_sram;
wire [0:1] mux_2level_tapbuf_size2_154_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_155_sram;
wire [0:1] mux_2level_tapbuf_size2_155_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_156_sram;
wire [0:1] mux_2level_tapbuf_size2_156_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_157_sram;
wire [0:1] mux_2level_tapbuf_size2_157_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_158_sram;
wire [0:1] mux_2level_tapbuf_size2_158_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_159_sram;
wire [0:1] mux_2level_tapbuf_size2_159_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_15_sram;
wire [0:1] mux_2level_tapbuf_size2_15_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_160_sram;
wire [0:1] mux_2level_tapbuf_size2_160_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_161_sram;
wire [0:1] mux_2level_tapbuf_size2_161_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_162_sram;
wire [0:1] mux_2level_tapbuf_size2_162_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_163_sram;
wire [0:1] mux_2level_tapbuf_size2_163_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_164_sram;
wire [0:1] mux_2level_tapbuf_size2_164_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_165_sram;
wire [0:1] mux_2level_tapbuf_size2_165_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_166_sram;
wire [0:1] mux_2level_tapbuf_size2_166_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_167_sram;
wire [0:1] mux_2level_tapbuf_size2_167_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_168_sram;
wire [0:1] mux_2level_tapbuf_size2_168_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_169_sram;
wire [0:1] mux_2level_tapbuf_size2_169_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_16_sram;
wire [0:1] mux_2level_tapbuf_size2_16_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_170_sram;
wire [0:1] mux_2level_tapbuf_size2_170_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_171_sram;
wire [0:1] mux_2level_tapbuf_size2_171_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_172_sram;
wire [0:1] mux_2level_tapbuf_size2_172_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_173_sram;
wire [0:1] mux_2level_tapbuf_size2_173_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_174_sram;
wire [0:1] mux_2level_tapbuf_size2_174_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_175_sram;
wire [0:1] mux_2level_tapbuf_size2_175_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_176_sram;
wire [0:1] mux_2level_tapbuf_size2_176_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_177_sram;
wire [0:1] mux_2level_tapbuf_size2_177_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_178_sram;
wire [0:1] mux_2level_tapbuf_size2_178_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_179_sram;
wire [0:1] mux_2level_tapbuf_size2_179_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_17_sram;
wire [0:1] mux_2level_tapbuf_size2_17_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_180_sram;
wire [0:1] mux_2level_tapbuf_size2_180_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_181_sram;
wire [0:1] mux_2level_tapbuf_size2_181_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_182_sram;
wire [0:1] mux_2level_tapbuf_size2_182_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_183_sram;
wire [0:1] mux_2level_tapbuf_size2_183_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_184_sram;
wire [0:1] mux_2level_tapbuf_size2_184_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_185_sram;
wire [0:1] mux_2level_tapbuf_size2_185_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_186_sram;
wire [0:1] mux_2level_tapbuf_size2_186_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_187_sram;
wire [0:1] mux_2level_tapbuf_size2_187_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_188_sram;
wire [0:1] mux_2level_tapbuf_size2_188_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_189_sram;
wire [0:1] mux_2level_tapbuf_size2_189_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_18_sram;
wire [0:1] mux_2level_tapbuf_size2_18_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_190_sram;
wire [0:1] mux_2level_tapbuf_size2_190_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_191_sram;
wire [0:1] mux_2level_tapbuf_size2_191_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_192_sram;
wire [0:1] mux_2level_tapbuf_size2_192_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_193_sram;
wire [0:1] mux_2level_tapbuf_size2_193_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_194_sram;
wire [0:1] mux_2level_tapbuf_size2_194_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_195_sram;
wire [0:1] mux_2level_tapbuf_size2_195_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_196_sram;
wire [0:1] mux_2level_tapbuf_size2_196_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_197_sram;
wire [0:1] mux_2level_tapbuf_size2_197_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_198_sram;
wire [0:1] mux_2level_tapbuf_size2_198_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_199_sram;
wire [0:1] mux_2level_tapbuf_size2_199_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_19_sram;
wire [0:1] mux_2level_tapbuf_size2_19_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_1_sram;
wire [0:1] mux_2level_tapbuf_size2_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_200_sram;
wire [0:1] mux_2level_tapbuf_size2_200_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_201_sram;
wire [0:1] mux_2level_tapbuf_size2_201_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_202_sram;
wire [0:1] mux_2level_tapbuf_size2_202_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_203_sram;
wire [0:1] mux_2level_tapbuf_size2_203_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_204_sram;
wire [0:1] mux_2level_tapbuf_size2_204_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_205_sram;
wire [0:1] mux_2level_tapbuf_size2_205_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_206_sram;
wire [0:1] mux_2level_tapbuf_size2_206_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_207_sram;
wire [0:1] mux_2level_tapbuf_size2_207_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_208_sram;
wire [0:1] mux_2level_tapbuf_size2_208_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_209_sram;
wire [0:1] mux_2level_tapbuf_size2_209_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_20_sram;
wire [0:1] mux_2level_tapbuf_size2_20_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_210_sram;
wire [0:1] mux_2level_tapbuf_size2_210_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_211_sram;
wire [0:1] mux_2level_tapbuf_size2_211_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_212_sram;
wire [0:1] mux_2level_tapbuf_size2_212_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_213_sram;
wire [0:1] mux_2level_tapbuf_size2_213_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_214_sram;
wire [0:1] mux_2level_tapbuf_size2_214_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_215_sram;
wire [0:1] mux_2level_tapbuf_size2_215_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_216_sram;
wire [0:1] mux_2level_tapbuf_size2_216_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_217_sram;
wire [0:1] mux_2level_tapbuf_size2_217_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_218_sram;
wire [0:1] mux_2level_tapbuf_size2_218_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_219_sram;
wire [0:1] mux_2level_tapbuf_size2_219_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_21_sram;
wire [0:1] mux_2level_tapbuf_size2_21_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_220_sram;
wire [0:1] mux_2level_tapbuf_size2_220_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_221_sram;
wire [0:1] mux_2level_tapbuf_size2_221_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_222_sram;
wire [0:1] mux_2level_tapbuf_size2_222_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_223_sram;
wire [0:1] mux_2level_tapbuf_size2_223_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_224_sram;
wire [0:1] mux_2level_tapbuf_size2_224_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_225_sram;
wire [0:1] mux_2level_tapbuf_size2_225_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_226_sram;
wire [0:1] mux_2level_tapbuf_size2_226_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_227_sram;
wire [0:1] mux_2level_tapbuf_size2_227_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_228_sram;
wire [0:1] mux_2level_tapbuf_size2_228_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_229_sram;
wire [0:1] mux_2level_tapbuf_size2_229_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_22_sram;
wire [0:1] mux_2level_tapbuf_size2_22_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_230_sram;
wire [0:1] mux_2level_tapbuf_size2_230_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_231_sram;
wire [0:1] mux_2level_tapbuf_size2_231_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_232_sram;
wire [0:1] mux_2level_tapbuf_size2_232_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_233_sram;
wire [0:1] mux_2level_tapbuf_size2_233_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_234_sram;
wire [0:1] mux_2level_tapbuf_size2_234_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_235_sram;
wire [0:1] mux_2level_tapbuf_size2_235_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_236_sram;
wire [0:1] mux_2level_tapbuf_size2_236_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_237_sram;
wire [0:1] mux_2level_tapbuf_size2_237_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_238_sram;
wire [0:1] mux_2level_tapbuf_size2_238_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_239_sram;
wire [0:1] mux_2level_tapbuf_size2_239_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_23_sram;
wire [0:1] mux_2level_tapbuf_size2_23_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_24_sram;
wire [0:1] mux_2level_tapbuf_size2_24_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_25_sram;
wire [0:1] mux_2level_tapbuf_size2_25_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_26_sram;
wire [0:1] mux_2level_tapbuf_size2_26_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_27_sram;
wire [0:1] mux_2level_tapbuf_size2_27_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_28_sram;
wire [0:1] mux_2level_tapbuf_size2_28_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_29_sram;
wire [0:1] mux_2level_tapbuf_size2_29_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_2_sram;
wire [0:1] mux_2level_tapbuf_size2_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_30_sram;
wire [0:1] mux_2level_tapbuf_size2_30_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_31_sram;
wire [0:1] mux_2level_tapbuf_size2_31_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_32_sram;
wire [0:1] mux_2level_tapbuf_size2_32_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_33_sram;
wire [0:1] mux_2level_tapbuf_size2_33_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_34_sram;
wire [0:1] mux_2level_tapbuf_size2_34_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_35_sram;
wire [0:1] mux_2level_tapbuf_size2_35_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_36_sram;
wire [0:1] mux_2level_tapbuf_size2_36_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_37_sram;
wire [0:1] mux_2level_tapbuf_size2_37_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_38_sram;
wire [0:1] mux_2level_tapbuf_size2_38_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_39_sram;
wire [0:1] mux_2level_tapbuf_size2_39_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_3_sram;
wire [0:1] mux_2level_tapbuf_size2_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_40_sram;
wire [0:1] mux_2level_tapbuf_size2_40_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_41_sram;
wire [0:1] mux_2level_tapbuf_size2_41_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_42_sram;
wire [0:1] mux_2level_tapbuf_size2_42_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_43_sram;
wire [0:1] mux_2level_tapbuf_size2_43_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_44_sram;
wire [0:1] mux_2level_tapbuf_size2_44_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_45_sram;
wire [0:1] mux_2level_tapbuf_size2_45_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_46_sram;
wire [0:1] mux_2level_tapbuf_size2_46_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_47_sram;
wire [0:1] mux_2level_tapbuf_size2_47_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_48_sram;
wire [0:1] mux_2level_tapbuf_size2_48_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_49_sram;
wire [0:1] mux_2level_tapbuf_size2_49_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_4_sram;
wire [0:1] mux_2level_tapbuf_size2_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_50_sram;
wire [0:1] mux_2level_tapbuf_size2_50_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_51_sram;
wire [0:1] mux_2level_tapbuf_size2_51_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_52_sram;
wire [0:1] mux_2level_tapbuf_size2_52_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_53_sram;
wire [0:1] mux_2level_tapbuf_size2_53_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_54_sram;
wire [0:1] mux_2level_tapbuf_size2_54_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_55_sram;
wire [0:1] mux_2level_tapbuf_size2_55_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_56_sram;
wire [0:1] mux_2level_tapbuf_size2_56_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_57_sram;
wire [0:1] mux_2level_tapbuf_size2_57_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_58_sram;
wire [0:1] mux_2level_tapbuf_size2_58_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_59_sram;
wire [0:1] mux_2level_tapbuf_size2_59_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_5_sram;
wire [0:1] mux_2level_tapbuf_size2_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_60_sram;
wire [0:1] mux_2level_tapbuf_size2_60_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_61_sram;
wire [0:1] mux_2level_tapbuf_size2_61_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_62_sram;
wire [0:1] mux_2level_tapbuf_size2_62_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_63_sram;
wire [0:1] mux_2level_tapbuf_size2_63_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_64_sram;
wire [0:1] mux_2level_tapbuf_size2_64_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_65_sram;
wire [0:1] mux_2level_tapbuf_size2_65_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_66_sram;
wire [0:1] mux_2level_tapbuf_size2_66_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_67_sram;
wire [0:1] mux_2level_tapbuf_size2_67_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_68_sram;
wire [0:1] mux_2level_tapbuf_size2_68_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_69_sram;
wire [0:1] mux_2level_tapbuf_size2_69_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_6_sram;
wire [0:1] mux_2level_tapbuf_size2_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_70_sram;
wire [0:1] mux_2level_tapbuf_size2_70_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_71_sram;
wire [0:1] mux_2level_tapbuf_size2_71_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_72_sram;
wire [0:1] mux_2level_tapbuf_size2_72_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_73_sram;
wire [0:1] mux_2level_tapbuf_size2_73_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_74_sram;
wire [0:1] mux_2level_tapbuf_size2_74_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_75_sram;
wire [0:1] mux_2level_tapbuf_size2_75_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_76_sram;
wire [0:1] mux_2level_tapbuf_size2_76_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_77_sram;
wire [0:1] mux_2level_tapbuf_size2_77_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_78_sram;
wire [0:1] mux_2level_tapbuf_size2_78_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_79_sram;
wire [0:1] mux_2level_tapbuf_size2_79_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_7_sram;
wire [0:1] mux_2level_tapbuf_size2_7_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_80_sram;
wire [0:1] mux_2level_tapbuf_size2_80_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_81_sram;
wire [0:1] mux_2level_tapbuf_size2_81_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_82_sram;
wire [0:1] mux_2level_tapbuf_size2_82_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_83_sram;
wire [0:1] mux_2level_tapbuf_size2_83_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_84_sram;
wire [0:1] mux_2level_tapbuf_size2_84_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_85_sram;
wire [0:1] mux_2level_tapbuf_size2_85_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_86_sram;
wire [0:1] mux_2level_tapbuf_size2_86_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_87_sram;
wire [0:1] mux_2level_tapbuf_size2_87_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_88_sram;
wire [0:1] mux_2level_tapbuf_size2_88_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_89_sram;
wire [0:1] mux_2level_tapbuf_size2_89_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_8_sram;
wire [0:1] mux_2level_tapbuf_size2_8_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_90_sram;
wire [0:1] mux_2level_tapbuf_size2_90_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_91_sram;
wire [0:1] mux_2level_tapbuf_size2_91_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_92_sram;
wire [0:1] mux_2level_tapbuf_size2_92_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_93_sram;
wire [0:1] mux_2level_tapbuf_size2_93_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_94_sram;
wire [0:1] mux_2level_tapbuf_size2_94_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_95_sram;
wire [0:1] mux_2level_tapbuf_size2_95_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_96_sram;
wire [0:1] mux_2level_tapbuf_size2_96_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_97_sram;
wire [0:1] mux_2level_tapbuf_size2_97_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_98_sram;
wire [0:1] mux_2level_tapbuf_size2_98_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_99_sram;
wire [0:1] mux_2level_tapbuf_size2_99_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_9_sram;
wire [0:1] mux_2level_tapbuf_size2_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_100_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_101_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_102_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_103_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_104_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_105_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_106_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_107_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_108_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_109_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_110_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_111_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_112_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_113_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_114_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_115_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_116_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_117_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_118_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_119_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_120_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_121_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_122_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_123_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_124_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_125_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_126_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_127_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_128_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_129_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_130_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_131_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_132_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_133_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_134_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_135_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_136_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_137_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_138_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_139_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_140_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_141_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_142_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_143_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_144_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_145_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_146_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_147_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_148_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_149_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_150_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_151_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_152_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_153_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_154_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_155_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_156_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_157_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_158_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_159_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_160_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_161_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_162_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_163_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_164_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_165_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_166_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_167_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_168_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_169_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_170_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_171_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_172_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_173_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_174_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_175_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_176_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_177_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_178_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_179_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_180_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_181_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_182_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_183_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_184_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_185_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_186_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_187_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_188_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_189_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_190_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_191_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_192_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_193_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_194_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_195_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_196_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_197_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_198_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_199_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_200_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_201_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_202_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_203_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_204_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_205_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_206_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_207_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_208_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_209_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_210_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_211_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_212_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_213_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_214_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_215_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_216_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_217_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_218_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_219_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_220_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_221_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_222_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_223_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_224_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_225_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_226_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_227_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_228_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_229_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_230_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_231_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_232_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_233_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_234_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_235_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_236_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_237_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_238_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_79_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_80_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_81_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_82_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_83_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_84_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_85_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_86_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_87_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_88_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_89_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_90_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_91_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_92_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_93_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_94_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_95_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_96_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_97_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_98_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_99_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[148] = chanx_right_in[0];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[139] = chanx_right_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[138] = chanx_right_in[10];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[129] = chanx_right_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[128] = chanx_right_in[20];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[119] = chanx_right_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[118] = chanx_right_in[30];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[109] = chanx_right_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[108] = chanx_right_in[40];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[99] = chanx_right_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[98] = chanx_right_in[50];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[89] = chanx_right_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[88] = chanx_right_in[60];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[79] = chanx_right_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[78] = chanx_right_in[70];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[69] = chanx_right_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[68] = chanx_right_in[80];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[59] = chanx_right_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[58] = chanx_right_in[90];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[49] = chanx_right_in[99];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[48] = chanx_right_in[100];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[39] = chanx_right_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[38] = chanx_right_in[110];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[29] = chanx_right_in[119];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[28] = chanx_right_in[120];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[19] = chanx_right_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[18] = chanx_right_in[130];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[9] = chanx_right_in[139];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[8] = chanx_right_in[140];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[149] = chanx_right_in[149];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[148] = chany_bottom_in[0];
// ----- Local connection due to Wire 167 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[139] = chany_bottom_in[9];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[138] = chany_bottom_in[10];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[129] = chany_bottom_in[19];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[128] = chany_bottom_in[20];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[119] = chany_bottom_in[29];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[118] = chany_bottom_in[30];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[109] = chany_bottom_in[39];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[108] = chany_bottom_in[40];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[99] = chany_bottom_in[49];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[98] = chany_bottom_in[50];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[89] = chany_bottom_in[59];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[88] = chany_bottom_in[60];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[79] = chany_bottom_in[69];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[78] = chany_bottom_in[70];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[69] = chany_bottom_in[79];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[68] = chany_bottom_in[80];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[59] = chany_bottom_in[89];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[58] = chany_bottom_in[90];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[49] = chany_bottom_in[99];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[48] = chany_bottom_in[100];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[39] = chany_bottom_in[109];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[38] = chany_bottom_in[110];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[29] = chany_bottom_in[119];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[28] = chany_bottom_in[120];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[19] = chany_bottom_in[129];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[18] = chany_bottom_in[130];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[9] = chany_bottom_in[139];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[8] = chany_bottom_in[140];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[149] = chany_bottom_in[149];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size2 mux_right_track_0 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[148]}),
		.sram(mux_2level_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_0_sram_inv[0:1]),
		.out(chanx_right_out[0]));

	mux_2level_tapbuf_size2 mux_right_track_2 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[147]}),
		.sram(mux_2level_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_1_sram_inv[0:1]),
		.out(chanx_right_out[1]));

	mux_2level_tapbuf_size2 mux_right_track_4 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[146]}),
		.sram(mux_2level_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_2_sram_inv[0:1]),
		.out(chanx_right_out[2]));

	mux_2level_tapbuf_size2 mux_right_track_6 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[145]}),
		.sram(mux_2level_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_3_sram_inv[0:1]),
		.out(chanx_right_out[3]));

	mux_2level_tapbuf_size2 mux_right_track_8 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[144]}),
		.sram(mux_2level_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_4_sram_inv[0:1]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size2 mux_right_track_10 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[143]}),
		.sram(mux_2level_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_5_sram_inv[0:1]),
		.out(chanx_right_out[5]));

	mux_2level_tapbuf_size2 mux_right_track_12 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[142]}),
		.sram(mux_2level_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_6_sram_inv[0:1]),
		.out(chanx_right_out[6]));

	mux_2level_tapbuf_size2 mux_right_track_14 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[141]}),
		.sram(mux_2level_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_7_sram_inv[0:1]),
		.out(chanx_right_out[7]));

	mux_2level_tapbuf_size2 mux_right_track_20 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[138]}),
		.sram(mux_2level_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_8_sram_inv[0:1]),
		.out(chanx_right_out[10]));

	mux_2level_tapbuf_size2 mux_right_track_22 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[137]}),
		.sram(mux_2level_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_9_sram_inv[0:1]),
		.out(chanx_right_out[11]));

	mux_2level_tapbuf_size2 mux_right_track_24 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[136]}),
		.sram(mux_2level_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_10_sram_inv[0:1]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size2 mux_right_track_26 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[135]}),
		.sram(mux_2level_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_11_sram_inv[0:1]),
		.out(chanx_right_out[13]));

	mux_2level_tapbuf_size2 mux_right_track_28 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[134]}),
		.sram(mux_2level_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_12_sram_inv[0:1]),
		.out(chanx_right_out[14]));

	mux_2level_tapbuf_size2 mux_right_track_30 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[133]}),
		.sram(mux_2level_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_13_sram_inv[0:1]),
		.out(chanx_right_out[15]));

	mux_2level_tapbuf_size2 mux_right_track_32 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[132]}),
		.sram(mux_2level_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_14_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size2 mux_right_track_34 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[131]}),
		.sram(mux_2level_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_15_sram_inv[0:1]),
		.out(chanx_right_out[17]));

	mux_2level_tapbuf_size2 mux_right_track_40 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[128]}),
		.sram(mux_2level_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_16_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size2 mux_right_track_42 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[127]}),
		.sram(mux_2level_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_17_sram_inv[0:1]),
		.out(chanx_right_out[21]));

	mux_2level_tapbuf_size2 mux_right_track_44 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[126]}),
		.sram(mux_2level_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_18_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_2level_tapbuf_size2 mux_right_track_46 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[125]}),
		.sram(mux_2level_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_19_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_2level_tapbuf_size2 mux_right_track_48 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[124]}),
		.sram(mux_2level_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_20_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size2 mux_right_track_50 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[123]}),
		.sram(mux_2level_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_21_sram_inv[0:1]),
		.out(chanx_right_out[25]));

	mux_2level_tapbuf_size2 mux_right_track_52 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[122]}),
		.sram(mux_2level_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_22_sram_inv[0:1]),
		.out(chanx_right_out[26]));

	mux_2level_tapbuf_size2 mux_right_track_54 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[121]}),
		.sram(mux_2level_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_23_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_2level_tapbuf_size2 mux_right_track_60 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[118]}),
		.sram(mux_2level_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_24_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_2level_tapbuf_size2 mux_right_track_62 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[117]}),
		.sram(mux_2level_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_25_sram_inv[0:1]),
		.out(chanx_right_out[31]));

	mux_2level_tapbuf_size2 mux_right_track_64 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[116]}),
		.sram(mux_2level_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_26_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size2 mux_right_track_66 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[115]}),
		.sram(mux_2level_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_27_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	mux_2level_tapbuf_size2 mux_right_track_68 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[114]}),
		.sram(mux_2level_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_28_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_2level_tapbuf_size2 mux_right_track_70 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[113]}),
		.sram(mux_2level_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_29_sram_inv[0:1]),
		.out(chanx_right_out[35]));

	mux_2level_tapbuf_size2 mux_right_track_72 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[112]}),
		.sram(mux_2level_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_30_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size2 mux_right_track_74 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[111]}),
		.sram(mux_2level_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_31_sram_inv[0:1]),
		.out(chanx_right_out[37]));

	mux_2level_tapbuf_size2 mux_right_track_80 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[108]}),
		.sram(mux_2level_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_32_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size2 mux_right_track_82 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[107]}),
		.sram(mux_2level_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_33_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	mux_2level_tapbuf_size2 mux_right_track_84 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[106]}),
		.sram(mux_2level_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_34_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_2level_tapbuf_size2 mux_right_track_86 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[105]}),
		.sram(mux_2level_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_35_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_2level_tapbuf_size2 mux_right_track_88 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[104]}),
		.sram(mux_2level_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_36_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	mux_2level_tapbuf_size2 mux_right_track_90 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[103]}),
		.sram(mux_2level_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_37_sram_inv[0:1]),
		.out(chanx_right_out[45]));

	mux_2level_tapbuf_size2 mux_right_track_92 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[102]}),
		.sram(mux_2level_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_38_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	mux_2level_tapbuf_size2 mux_right_track_94 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[101]}),
		.sram(mux_2level_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_39_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_2level_tapbuf_size2 mux_right_track_100 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[98]}),
		.sram(mux_2level_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_40_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	mux_2level_tapbuf_size2 mux_right_track_102 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[97]}),
		.sram(mux_2level_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_41_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	mux_2level_tapbuf_size2 mux_right_track_104 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[96]}),
		.sram(mux_2level_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_42_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	mux_2level_tapbuf_size2 mux_right_track_106 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[95]}),
		.sram(mux_2level_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_43_sram_inv[0:1]),
		.out(chanx_right_out[53]));

	mux_2level_tapbuf_size2 mux_right_track_108 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[94]}),
		.sram(mux_2level_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_44_sram_inv[0:1]),
		.out(chanx_right_out[54]));

	mux_2level_tapbuf_size2 mux_right_track_110 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[93]}),
		.sram(mux_2level_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_45_sram_inv[0:1]),
		.out(chanx_right_out[55]));

	mux_2level_tapbuf_size2 mux_right_track_112 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[92]}),
		.sram(mux_2level_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_46_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_2level_tapbuf_size2 mux_right_track_114 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[91]}),
		.sram(mux_2level_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_47_sram_inv[0:1]),
		.out(chanx_right_out[57]));

	mux_2level_tapbuf_size2 mux_right_track_120 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[88]}),
		.sram(mux_2level_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_48_sram_inv[0:1]),
		.out(chanx_right_out[60]));

	mux_2level_tapbuf_size2 mux_right_track_122 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[87]}),
		.sram(mux_2level_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_49_sram_inv[0:1]),
		.out(chanx_right_out[61]));

	mux_2level_tapbuf_size2 mux_right_track_124 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[86]}),
		.sram(mux_2level_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_50_sram_inv[0:1]),
		.out(chanx_right_out[62]));

	mux_2level_tapbuf_size2 mux_right_track_126 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[85]}),
		.sram(mux_2level_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_51_sram_inv[0:1]),
		.out(chanx_right_out[63]));

	mux_2level_tapbuf_size2 mux_right_track_128 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[84]}),
		.sram(mux_2level_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_52_sram_inv[0:1]),
		.out(chanx_right_out[64]));

	mux_2level_tapbuf_size2 mux_right_track_130 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[83]}),
		.sram(mux_2level_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_53_sram_inv[0:1]),
		.out(chanx_right_out[65]));

	mux_2level_tapbuf_size2 mux_right_track_132 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[82]}),
		.sram(mux_2level_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_54_sram_inv[0:1]),
		.out(chanx_right_out[66]));

	mux_2level_tapbuf_size2 mux_right_track_134 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[81]}),
		.sram(mux_2level_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_55_sram_inv[0:1]),
		.out(chanx_right_out[67]));

	mux_2level_tapbuf_size2 mux_right_track_140 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[78]}),
		.sram(mux_2level_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_56_sram_inv[0:1]),
		.out(chanx_right_out[70]));

	mux_2level_tapbuf_size2 mux_right_track_142 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[77]}),
		.sram(mux_2level_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_57_sram_inv[0:1]),
		.out(chanx_right_out[71]));

	mux_2level_tapbuf_size2 mux_right_track_144 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[76]}),
		.sram(mux_2level_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_58_sram_inv[0:1]),
		.out(chanx_right_out[72]));

	mux_2level_tapbuf_size2 mux_right_track_146 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[75]}),
		.sram(mux_2level_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_59_sram_inv[0:1]),
		.out(chanx_right_out[73]));

	mux_2level_tapbuf_size2 mux_right_track_148 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[74]}),
		.sram(mux_2level_tapbuf_size2_60_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_60_sram_inv[0:1]),
		.out(chanx_right_out[74]));

	mux_2level_tapbuf_size2 mux_right_track_150 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[73]}),
		.sram(mux_2level_tapbuf_size2_61_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_61_sram_inv[0:1]),
		.out(chanx_right_out[75]));

	mux_2level_tapbuf_size2 mux_right_track_152 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[72]}),
		.sram(mux_2level_tapbuf_size2_62_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_62_sram_inv[0:1]),
		.out(chanx_right_out[76]));

	mux_2level_tapbuf_size2 mux_right_track_154 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[71]}),
		.sram(mux_2level_tapbuf_size2_63_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_63_sram_inv[0:1]),
		.out(chanx_right_out[77]));

	mux_2level_tapbuf_size2 mux_right_track_160 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[68]}),
		.sram(mux_2level_tapbuf_size2_64_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_64_sram_inv[0:1]),
		.out(chanx_right_out[80]));

	mux_2level_tapbuf_size2 mux_right_track_162 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[67]}),
		.sram(mux_2level_tapbuf_size2_65_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_65_sram_inv[0:1]),
		.out(chanx_right_out[81]));

	mux_2level_tapbuf_size2 mux_right_track_164 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[66]}),
		.sram(mux_2level_tapbuf_size2_66_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_66_sram_inv[0:1]),
		.out(chanx_right_out[82]));

	mux_2level_tapbuf_size2 mux_right_track_166 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[65]}),
		.sram(mux_2level_tapbuf_size2_67_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_67_sram_inv[0:1]),
		.out(chanx_right_out[83]));

	mux_2level_tapbuf_size2 mux_right_track_168 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[64]}),
		.sram(mux_2level_tapbuf_size2_68_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_68_sram_inv[0:1]),
		.out(chanx_right_out[84]));

	mux_2level_tapbuf_size2 mux_right_track_170 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[63]}),
		.sram(mux_2level_tapbuf_size2_69_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_69_sram_inv[0:1]),
		.out(chanx_right_out[85]));

	mux_2level_tapbuf_size2 mux_right_track_172 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[62]}),
		.sram(mux_2level_tapbuf_size2_70_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_70_sram_inv[0:1]),
		.out(chanx_right_out[86]));

	mux_2level_tapbuf_size2 mux_right_track_174 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[61]}),
		.sram(mux_2level_tapbuf_size2_71_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_71_sram_inv[0:1]),
		.out(chanx_right_out[87]));

	mux_2level_tapbuf_size2 mux_right_track_180 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[58]}),
		.sram(mux_2level_tapbuf_size2_72_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_72_sram_inv[0:1]),
		.out(chanx_right_out[90]));

	mux_2level_tapbuf_size2 mux_right_track_182 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[57]}),
		.sram(mux_2level_tapbuf_size2_73_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_73_sram_inv[0:1]),
		.out(chanx_right_out[91]));

	mux_2level_tapbuf_size2 mux_right_track_184 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[56]}),
		.sram(mux_2level_tapbuf_size2_74_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_74_sram_inv[0:1]),
		.out(chanx_right_out[92]));

	mux_2level_tapbuf_size2 mux_right_track_186 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[55]}),
		.sram(mux_2level_tapbuf_size2_75_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_75_sram_inv[0:1]),
		.out(chanx_right_out[93]));

	mux_2level_tapbuf_size2 mux_right_track_188 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[54]}),
		.sram(mux_2level_tapbuf_size2_76_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_76_sram_inv[0:1]),
		.out(chanx_right_out[94]));

	mux_2level_tapbuf_size2 mux_right_track_190 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[53]}),
		.sram(mux_2level_tapbuf_size2_77_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_77_sram_inv[0:1]),
		.out(chanx_right_out[95]));

	mux_2level_tapbuf_size2 mux_right_track_192 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[52]}),
		.sram(mux_2level_tapbuf_size2_78_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_78_sram_inv[0:1]),
		.out(chanx_right_out[96]));

	mux_2level_tapbuf_size2 mux_right_track_194 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[51]}),
		.sram(mux_2level_tapbuf_size2_79_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_79_sram_inv[0:1]),
		.out(chanx_right_out[97]));

	mux_2level_tapbuf_size2 mux_right_track_200 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[48]}),
		.sram(mux_2level_tapbuf_size2_80_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_80_sram_inv[0:1]),
		.out(chanx_right_out[100]));

	mux_2level_tapbuf_size2 mux_right_track_202 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[47]}),
		.sram(mux_2level_tapbuf_size2_81_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_81_sram_inv[0:1]),
		.out(chanx_right_out[101]));

	mux_2level_tapbuf_size2 mux_right_track_204 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[46]}),
		.sram(mux_2level_tapbuf_size2_82_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_82_sram_inv[0:1]),
		.out(chanx_right_out[102]));

	mux_2level_tapbuf_size2 mux_right_track_206 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[45]}),
		.sram(mux_2level_tapbuf_size2_83_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_83_sram_inv[0:1]),
		.out(chanx_right_out[103]));

	mux_2level_tapbuf_size2 mux_right_track_208 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[44]}),
		.sram(mux_2level_tapbuf_size2_84_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_84_sram_inv[0:1]),
		.out(chanx_right_out[104]));

	mux_2level_tapbuf_size2 mux_right_track_210 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[43]}),
		.sram(mux_2level_tapbuf_size2_85_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_85_sram_inv[0:1]),
		.out(chanx_right_out[105]));

	mux_2level_tapbuf_size2 mux_right_track_212 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[42]}),
		.sram(mux_2level_tapbuf_size2_86_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_86_sram_inv[0:1]),
		.out(chanx_right_out[106]));

	mux_2level_tapbuf_size2 mux_right_track_214 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[41]}),
		.sram(mux_2level_tapbuf_size2_87_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_87_sram_inv[0:1]),
		.out(chanx_right_out[107]));

	mux_2level_tapbuf_size2 mux_right_track_220 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[38]}),
		.sram(mux_2level_tapbuf_size2_88_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_88_sram_inv[0:1]),
		.out(chanx_right_out[110]));

	mux_2level_tapbuf_size2 mux_right_track_222 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[37]}),
		.sram(mux_2level_tapbuf_size2_89_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_89_sram_inv[0:1]),
		.out(chanx_right_out[111]));

	mux_2level_tapbuf_size2 mux_right_track_224 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[36]}),
		.sram(mux_2level_tapbuf_size2_90_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_90_sram_inv[0:1]),
		.out(chanx_right_out[112]));

	mux_2level_tapbuf_size2 mux_right_track_226 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[35]}),
		.sram(mux_2level_tapbuf_size2_91_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_91_sram_inv[0:1]),
		.out(chanx_right_out[113]));

	mux_2level_tapbuf_size2 mux_right_track_228 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[34]}),
		.sram(mux_2level_tapbuf_size2_92_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_92_sram_inv[0:1]),
		.out(chanx_right_out[114]));

	mux_2level_tapbuf_size2 mux_right_track_230 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[33]}),
		.sram(mux_2level_tapbuf_size2_93_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_93_sram_inv[0:1]),
		.out(chanx_right_out[115]));

	mux_2level_tapbuf_size2 mux_right_track_232 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[32]}),
		.sram(mux_2level_tapbuf_size2_94_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_94_sram_inv[0:1]),
		.out(chanx_right_out[116]));

	mux_2level_tapbuf_size2 mux_right_track_234 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[31]}),
		.sram(mux_2level_tapbuf_size2_95_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_95_sram_inv[0:1]),
		.out(chanx_right_out[117]));

	mux_2level_tapbuf_size2 mux_right_track_240 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[28]}),
		.sram(mux_2level_tapbuf_size2_96_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_96_sram_inv[0:1]),
		.out(chanx_right_out[120]));

	mux_2level_tapbuf_size2 mux_right_track_242 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[27]}),
		.sram(mux_2level_tapbuf_size2_97_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_97_sram_inv[0:1]),
		.out(chanx_right_out[121]));

	mux_2level_tapbuf_size2 mux_right_track_244 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[26]}),
		.sram(mux_2level_tapbuf_size2_98_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_98_sram_inv[0:1]),
		.out(chanx_right_out[122]));

	mux_2level_tapbuf_size2 mux_right_track_246 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[25]}),
		.sram(mux_2level_tapbuf_size2_99_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_99_sram_inv[0:1]),
		.out(chanx_right_out[123]));

	mux_2level_tapbuf_size2 mux_right_track_248 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[24]}),
		.sram(mux_2level_tapbuf_size2_100_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_100_sram_inv[0:1]),
		.out(chanx_right_out[124]));

	mux_2level_tapbuf_size2 mux_right_track_250 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[23]}),
		.sram(mux_2level_tapbuf_size2_101_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_101_sram_inv[0:1]),
		.out(chanx_right_out[125]));

	mux_2level_tapbuf_size2 mux_right_track_252 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[22]}),
		.sram(mux_2level_tapbuf_size2_102_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_102_sram_inv[0:1]),
		.out(chanx_right_out[126]));

	mux_2level_tapbuf_size2 mux_right_track_254 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[21]}),
		.sram(mux_2level_tapbuf_size2_103_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_103_sram_inv[0:1]),
		.out(chanx_right_out[127]));

	mux_2level_tapbuf_size2 mux_right_track_260 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[18]}),
		.sram(mux_2level_tapbuf_size2_104_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_104_sram_inv[0:1]),
		.out(chanx_right_out[130]));

	mux_2level_tapbuf_size2 mux_right_track_262 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[17]}),
		.sram(mux_2level_tapbuf_size2_105_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_105_sram_inv[0:1]),
		.out(chanx_right_out[131]));

	mux_2level_tapbuf_size2 mux_right_track_264 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[16]}),
		.sram(mux_2level_tapbuf_size2_106_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_106_sram_inv[0:1]),
		.out(chanx_right_out[132]));

	mux_2level_tapbuf_size2 mux_right_track_266 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[15]}),
		.sram(mux_2level_tapbuf_size2_107_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_107_sram_inv[0:1]),
		.out(chanx_right_out[133]));

	mux_2level_tapbuf_size2 mux_right_track_268 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[14]}),
		.sram(mux_2level_tapbuf_size2_108_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_108_sram_inv[0:1]),
		.out(chanx_right_out[134]));

	mux_2level_tapbuf_size2 mux_right_track_270 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[13]}),
		.sram(mux_2level_tapbuf_size2_109_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_109_sram_inv[0:1]),
		.out(chanx_right_out[135]));

	mux_2level_tapbuf_size2 mux_right_track_272 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[12]}),
		.sram(mux_2level_tapbuf_size2_110_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_110_sram_inv[0:1]),
		.out(chanx_right_out[136]));

	mux_2level_tapbuf_size2 mux_right_track_274 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[11]}),
		.sram(mux_2level_tapbuf_size2_111_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_111_sram_inv[0:1]),
		.out(chanx_right_out[137]));

	mux_2level_tapbuf_size2 mux_right_track_280 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[8]}),
		.sram(mux_2level_tapbuf_size2_112_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_112_sram_inv[0:1]),
		.out(chanx_right_out[140]));

	mux_2level_tapbuf_size2 mux_right_track_282 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[7]}),
		.sram(mux_2level_tapbuf_size2_113_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_113_sram_inv[0:1]),
		.out(chanx_right_out[141]));

	mux_2level_tapbuf_size2 mux_right_track_284 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[6]}),
		.sram(mux_2level_tapbuf_size2_114_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_114_sram_inv[0:1]),
		.out(chanx_right_out[142]));

	mux_2level_tapbuf_size2 mux_right_track_286 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[5]}),
		.sram(mux_2level_tapbuf_size2_115_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_115_sram_inv[0:1]),
		.out(chanx_right_out[143]));

	mux_2level_tapbuf_size2 mux_right_track_288 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[4]}),
		.sram(mux_2level_tapbuf_size2_116_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_116_sram_inv[0:1]),
		.out(chanx_right_out[144]));

	mux_2level_tapbuf_size2 mux_right_track_290 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[3]}),
		.sram(mux_2level_tapbuf_size2_117_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_117_sram_inv[0:1]),
		.out(chanx_right_out[145]));

	mux_2level_tapbuf_size2 mux_right_track_292 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[2]}),
		.sram(mux_2level_tapbuf_size2_118_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_118_sram_inv[0:1]),
		.out(chanx_right_out[146]));

	mux_2level_tapbuf_size2 mux_right_track_294 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[1]}),
		.sram(mux_2level_tapbuf_size2_119_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_119_sram_inv[0:1]),
		.out(chanx_right_out[147]));

	mux_2level_tapbuf_size2 mux_bottom_track_1 (
		.in({chanx_right_in[148], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_120_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_120_sram_inv[0:1]),
		.out(chany_bottom_out[0]));

	mux_2level_tapbuf_size2 mux_bottom_track_3 (
		.in({chanx_right_in[147], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_121_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_121_sram_inv[0:1]),
		.out(chany_bottom_out[1]));

	mux_2level_tapbuf_size2 mux_bottom_track_5 (
		.in({chanx_right_in[146], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_122_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_122_sram_inv[0:1]),
		.out(chany_bottom_out[2]));

	mux_2level_tapbuf_size2 mux_bottom_track_7 (
		.in({chanx_right_in[145], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_123_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_123_sram_inv[0:1]),
		.out(chany_bottom_out[3]));

	mux_2level_tapbuf_size2 mux_bottom_track_9 (
		.in({chanx_right_in[144], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_124_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_124_sram_inv[0:1]),
		.out(chany_bottom_out[4]));

	mux_2level_tapbuf_size2 mux_bottom_track_11 (
		.in({chanx_right_in[143], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_125_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_125_sram_inv[0:1]),
		.out(chany_bottom_out[5]));

	mux_2level_tapbuf_size2 mux_bottom_track_13 (
		.in({chanx_right_in[142], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_126_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_126_sram_inv[0:1]),
		.out(chany_bottom_out[6]));

	mux_2level_tapbuf_size2 mux_bottom_track_15 (
		.in({chanx_right_in[141], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_127_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_127_sram_inv[0:1]),
		.out(chany_bottom_out[7]));

	mux_2level_tapbuf_size2 mux_bottom_track_21 (
		.in({chanx_right_in[138], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_128_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_128_sram_inv[0:1]),
		.out(chany_bottom_out[10]));

	mux_2level_tapbuf_size2 mux_bottom_track_23 (
		.in({chanx_right_in[137], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_129_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_129_sram_inv[0:1]),
		.out(chany_bottom_out[11]));

	mux_2level_tapbuf_size2 mux_bottom_track_25 (
		.in({chanx_right_in[136], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_130_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_130_sram_inv[0:1]),
		.out(chany_bottom_out[12]));

	mux_2level_tapbuf_size2 mux_bottom_track_27 (
		.in({chanx_right_in[135], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_131_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_131_sram_inv[0:1]),
		.out(chany_bottom_out[13]));

	mux_2level_tapbuf_size2 mux_bottom_track_29 (
		.in({chanx_right_in[134], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_132_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_132_sram_inv[0:1]),
		.out(chany_bottom_out[14]));

	mux_2level_tapbuf_size2 mux_bottom_track_31 (
		.in({chanx_right_in[133], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_133_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_133_sram_inv[0:1]),
		.out(chany_bottom_out[15]));

	mux_2level_tapbuf_size2 mux_bottom_track_33 (
		.in({chanx_right_in[132], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_134_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_134_sram_inv[0:1]),
		.out(chany_bottom_out[16]));

	mux_2level_tapbuf_size2 mux_bottom_track_35 (
		.in({chanx_right_in[131], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_135_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_135_sram_inv[0:1]),
		.out(chany_bottom_out[17]));

	mux_2level_tapbuf_size2 mux_bottom_track_41 (
		.in({chanx_right_in[128], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_136_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_136_sram_inv[0:1]),
		.out(chany_bottom_out[20]));

	mux_2level_tapbuf_size2 mux_bottom_track_43 (
		.in({chanx_right_in[127], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_137_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_137_sram_inv[0:1]),
		.out(chany_bottom_out[21]));

	mux_2level_tapbuf_size2 mux_bottom_track_45 (
		.in({chanx_right_in[126], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_138_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_138_sram_inv[0:1]),
		.out(chany_bottom_out[22]));

	mux_2level_tapbuf_size2 mux_bottom_track_47 (
		.in({chanx_right_in[125], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_139_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_139_sram_inv[0:1]),
		.out(chany_bottom_out[23]));

	mux_2level_tapbuf_size2 mux_bottom_track_49 (
		.in({chanx_right_in[124], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_140_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_140_sram_inv[0:1]),
		.out(chany_bottom_out[24]));

	mux_2level_tapbuf_size2 mux_bottom_track_51 (
		.in({chanx_right_in[123], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_141_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_141_sram_inv[0:1]),
		.out(chany_bottom_out[25]));

	mux_2level_tapbuf_size2 mux_bottom_track_53 (
		.in({chanx_right_in[122], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_142_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_142_sram_inv[0:1]),
		.out(chany_bottom_out[26]));

	mux_2level_tapbuf_size2 mux_bottom_track_55 (
		.in({chanx_right_in[121], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_143_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_143_sram_inv[0:1]),
		.out(chany_bottom_out[27]));

	mux_2level_tapbuf_size2 mux_bottom_track_61 (
		.in({chanx_right_in[118], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_144_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_144_sram_inv[0:1]),
		.out(chany_bottom_out[30]));

	mux_2level_tapbuf_size2 mux_bottom_track_63 (
		.in({chanx_right_in[117], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_145_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_145_sram_inv[0:1]),
		.out(chany_bottom_out[31]));

	mux_2level_tapbuf_size2 mux_bottom_track_65 (
		.in({chanx_right_in[116], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_146_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_146_sram_inv[0:1]),
		.out(chany_bottom_out[32]));

	mux_2level_tapbuf_size2 mux_bottom_track_67 (
		.in({chanx_right_in[115], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_147_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_147_sram_inv[0:1]),
		.out(chany_bottom_out[33]));

	mux_2level_tapbuf_size2 mux_bottom_track_69 (
		.in({chanx_right_in[114], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_148_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_148_sram_inv[0:1]),
		.out(chany_bottom_out[34]));

	mux_2level_tapbuf_size2 mux_bottom_track_71 (
		.in({chanx_right_in[113], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_149_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_149_sram_inv[0:1]),
		.out(chany_bottom_out[35]));

	mux_2level_tapbuf_size2 mux_bottom_track_73 (
		.in({chanx_right_in[112], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_150_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_150_sram_inv[0:1]),
		.out(chany_bottom_out[36]));

	mux_2level_tapbuf_size2 mux_bottom_track_75 (
		.in({chanx_right_in[111], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_151_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_151_sram_inv[0:1]),
		.out(chany_bottom_out[37]));

	mux_2level_tapbuf_size2 mux_bottom_track_81 (
		.in({chanx_right_in[108], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_152_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_152_sram_inv[0:1]),
		.out(chany_bottom_out[40]));

	mux_2level_tapbuf_size2 mux_bottom_track_83 (
		.in({chanx_right_in[107], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_153_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_153_sram_inv[0:1]),
		.out(chany_bottom_out[41]));

	mux_2level_tapbuf_size2 mux_bottom_track_85 (
		.in({chanx_right_in[106], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_154_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_154_sram_inv[0:1]),
		.out(chany_bottom_out[42]));

	mux_2level_tapbuf_size2 mux_bottom_track_87 (
		.in({chanx_right_in[105], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_155_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_155_sram_inv[0:1]),
		.out(chany_bottom_out[43]));

	mux_2level_tapbuf_size2 mux_bottom_track_89 (
		.in({chanx_right_in[104], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_156_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_156_sram_inv[0:1]),
		.out(chany_bottom_out[44]));

	mux_2level_tapbuf_size2 mux_bottom_track_91 (
		.in({chanx_right_in[103], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_157_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_157_sram_inv[0:1]),
		.out(chany_bottom_out[45]));

	mux_2level_tapbuf_size2 mux_bottom_track_93 (
		.in({chanx_right_in[102], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_158_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_158_sram_inv[0:1]),
		.out(chany_bottom_out[46]));

	mux_2level_tapbuf_size2 mux_bottom_track_95 (
		.in({chanx_right_in[101], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_159_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_159_sram_inv[0:1]),
		.out(chany_bottom_out[47]));

	mux_2level_tapbuf_size2 mux_bottom_track_101 (
		.in({chanx_right_in[98], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_160_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_160_sram_inv[0:1]),
		.out(chany_bottom_out[50]));

	mux_2level_tapbuf_size2 mux_bottom_track_103 (
		.in({chanx_right_in[97], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_161_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_161_sram_inv[0:1]),
		.out(chany_bottom_out[51]));

	mux_2level_tapbuf_size2 mux_bottom_track_105 (
		.in({chanx_right_in[96], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_162_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_162_sram_inv[0:1]),
		.out(chany_bottom_out[52]));

	mux_2level_tapbuf_size2 mux_bottom_track_107 (
		.in({chanx_right_in[95], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_163_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_163_sram_inv[0:1]),
		.out(chany_bottom_out[53]));

	mux_2level_tapbuf_size2 mux_bottom_track_109 (
		.in({chanx_right_in[94], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_164_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_164_sram_inv[0:1]),
		.out(chany_bottom_out[54]));

	mux_2level_tapbuf_size2 mux_bottom_track_111 (
		.in({chanx_right_in[93], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_165_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_165_sram_inv[0:1]),
		.out(chany_bottom_out[55]));

	mux_2level_tapbuf_size2 mux_bottom_track_113 (
		.in({chanx_right_in[92], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_166_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_166_sram_inv[0:1]),
		.out(chany_bottom_out[56]));

	mux_2level_tapbuf_size2 mux_bottom_track_115 (
		.in({chanx_right_in[91], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_167_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_167_sram_inv[0:1]),
		.out(chany_bottom_out[57]));

	mux_2level_tapbuf_size2 mux_bottom_track_121 (
		.in({chanx_right_in[88], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_168_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_168_sram_inv[0:1]),
		.out(chany_bottom_out[60]));

	mux_2level_tapbuf_size2 mux_bottom_track_123 (
		.in({chanx_right_in[87], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_169_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_169_sram_inv[0:1]),
		.out(chany_bottom_out[61]));

	mux_2level_tapbuf_size2 mux_bottom_track_125 (
		.in({chanx_right_in[86], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_170_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_170_sram_inv[0:1]),
		.out(chany_bottom_out[62]));

	mux_2level_tapbuf_size2 mux_bottom_track_127 (
		.in({chanx_right_in[85], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_171_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_171_sram_inv[0:1]),
		.out(chany_bottom_out[63]));

	mux_2level_tapbuf_size2 mux_bottom_track_129 (
		.in({chanx_right_in[84], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_172_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_172_sram_inv[0:1]),
		.out(chany_bottom_out[64]));

	mux_2level_tapbuf_size2 mux_bottom_track_131 (
		.in({chanx_right_in[83], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_173_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_173_sram_inv[0:1]),
		.out(chany_bottom_out[65]));

	mux_2level_tapbuf_size2 mux_bottom_track_133 (
		.in({chanx_right_in[82], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_174_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_174_sram_inv[0:1]),
		.out(chany_bottom_out[66]));

	mux_2level_tapbuf_size2 mux_bottom_track_135 (
		.in({chanx_right_in[81], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_175_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_175_sram_inv[0:1]),
		.out(chany_bottom_out[67]));

	mux_2level_tapbuf_size2 mux_bottom_track_141 (
		.in({chanx_right_in[78], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_176_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_176_sram_inv[0:1]),
		.out(chany_bottom_out[70]));

	mux_2level_tapbuf_size2 mux_bottom_track_143 (
		.in({chanx_right_in[77], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_177_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_177_sram_inv[0:1]),
		.out(chany_bottom_out[71]));

	mux_2level_tapbuf_size2 mux_bottom_track_145 (
		.in({chanx_right_in[76], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_178_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_178_sram_inv[0:1]),
		.out(chany_bottom_out[72]));

	mux_2level_tapbuf_size2 mux_bottom_track_147 (
		.in({chanx_right_in[75], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_179_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_179_sram_inv[0:1]),
		.out(chany_bottom_out[73]));

	mux_2level_tapbuf_size2 mux_bottom_track_149 (
		.in({chanx_right_in[74], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_180_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_180_sram_inv[0:1]),
		.out(chany_bottom_out[74]));

	mux_2level_tapbuf_size2 mux_bottom_track_151 (
		.in({chanx_right_in[73], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_181_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_181_sram_inv[0:1]),
		.out(chany_bottom_out[75]));

	mux_2level_tapbuf_size2 mux_bottom_track_153 (
		.in({chanx_right_in[72], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_182_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_182_sram_inv[0:1]),
		.out(chany_bottom_out[76]));

	mux_2level_tapbuf_size2 mux_bottom_track_155 (
		.in({chanx_right_in[71], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_183_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_183_sram_inv[0:1]),
		.out(chany_bottom_out[77]));

	mux_2level_tapbuf_size2 mux_bottom_track_161 (
		.in({chanx_right_in[68], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_184_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_184_sram_inv[0:1]),
		.out(chany_bottom_out[80]));

	mux_2level_tapbuf_size2 mux_bottom_track_163 (
		.in({chanx_right_in[67], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_185_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_185_sram_inv[0:1]),
		.out(chany_bottom_out[81]));

	mux_2level_tapbuf_size2 mux_bottom_track_165 (
		.in({chanx_right_in[66], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_186_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_186_sram_inv[0:1]),
		.out(chany_bottom_out[82]));

	mux_2level_tapbuf_size2 mux_bottom_track_167 (
		.in({chanx_right_in[65], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_187_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_187_sram_inv[0:1]),
		.out(chany_bottom_out[83]));

	mux_2level_tapbuf_size2 mux_bottom_track_169 (
		.in({chanx_right_in[64], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_188_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_188_sram_inv[0:1]),
		.out(chany_bottom_out[84]));

	mux_2level_tapbuf_size2 mux_bottom_track_171 (
		.in({chanx_right_in[63], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_189_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_189_sram_inv[0:1]),
		.out(chany_bottom_out[85]));

	mux_2level_tapbuf_size2 mux_bottom_track_173 (
		.in({chanx_right_in[62], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_190_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_190_sram_inv[0:1]),
		.out(chany_bottom_out[86]));

	mux_2level_tapbuf_size2 mux_bottom_track_175 (
		.in({chanx_right_in[61], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_191_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_191_sram_inv[0:1]),
		.out(chany_bottom_out[87]));

	mux_2level_tapbuf_size2 mux_bottom_track_181 (
		.in({chanx_right_in[58], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_192_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_192_sram_inv[0:1]),
		.out(chany_bottom_out[90]));

	mux_2level_tapbuf_size2 mux_bottom_track_183 (
		.in({chanx_right_in[57], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_193_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_193_sram_inv[0:1]),
		.out(chany_bottom_out[91]));

	mux_2level_tapbuf_size2 mux_bottom_track_185 (
		.in({chanx_right_in[56], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_194_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_194_sram_inv[0:1]),
		.out(chany_bottom_out[92]));

	mux_2level_tapbuf_size2 mux_bottom_track_187 (
		.in({chanx_right_in[55], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_195_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_195_sram_inv[0:1]),
		.out(chany_bottom_out[93]));

	mux_2level_tapbuf_size2 mux_bottom_track_189 (
		.in({chanx_right_in[54], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_196_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_196_sram_inv[0:1]),
		.out(chany_bottom_out[94]));

	mux_2level_tapbuf_size2 mux_bottom_track_191 (
		.in({chanx_right_in[53], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_197_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_197_sram_inv[0:1]),
		.out(chany_bottom_out[95]));

	mux_2level_tapbuf_size2 mux_bottom_track_193 (
		.in({chanx_right_in[52], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_198_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_198_sram_inv[0:1]),
		.out(chany_bottom_out[96]));

	mux_2level_tapbuf_size2 mux_bottom_track_195 (
		.in({chanx_right_in[51], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_199_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_199_sram_inv[0:1]),
		.out(chany_bottom_out[97]));

	mux_2level_tapbuf_size2 mux_bottom_track_201 (
		.in({chanx_right_in[48], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_200_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_200_sram_inv[0:1]),
		.out(chany_bottom_out[100]));

	mux_2level_tapbuf_size2 mux_bottom_track_203 (
		.in({chanx_right_in[47], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_201_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_201_sram_inv[0:1]),
		.out(chany_bottom_out[101]));

	mux_2level_tapbuf_size2 mux_bottom_track_205 (
		.in({chanx_right_in[46], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_202_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_202_sram_inv[0:1]),
		.out(chany_bottom_out[102]));

	mux_2level_tapbuf_size2 mux_bottom_track_207 (
		.in({chanx_right_in[45], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_203_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_203_sram_inv[0:1]),
		.out(chany_bottom_out[103]));

	mux_2level_tapbuf_size2 mux_bottom_track_209 (
		.in({chanx_right_in[44], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_204_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_204_sram_inv[0:1]),
		.out(chany_bottom_out[104]));

	mux_2level_tapbuf_size2 mux_bottom_track_211 (
		.in({chanx_right_in[43], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_205_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_205_sram_inv[0:1]),
		.out(chany_bottom_out[105]));

	mux_2level_tapbuf_size2 mux_bottom_track_213 (
		.in({chanx_right_in[42], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_206_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_206_sram_inv[0:1]),
		.out(chany_bottom_out[106]));

	mux_2level_tapbuf_size2 mux_bottom_track_215 (
		.in({chanx_right_in[41], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_207_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_207_sram_inv[0:1]),
		.out(chany_bottom_out[107]));

	mux_2level_tapbuf_size2 mux_bottom_track_221 (
		.in({chanx_right_in[38], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_208_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_208_sram_inv[0:1]),
		.out(chany_bottom_out[110]));

	mux_2level_tapbuf_size2 mux_bottom_track_223 (
		.in({chanx_right_in[37], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_209_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_209_sram_inv[0:1]),
		.out(chany_bottom_out[111]));

	mux_2level_tapbuf_size2 mux_bottom_track_225 (
		.in({chanx_right_in[36], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_210_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_210_sram_inv[0:1]),
		.out(chany_bottom_out[112]));

	mux_2level_tapbuf_size2 mux_bottom_track_227 (
		.in({chanx_right_in[35], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_211_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_211_sram_inv[0:1]),
		.out(chany_bottom_out[113]));

	mux_2level_tapbuf_size2 mux_bottom_track_229 (
		.in({chanx_right_in[34], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_212_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_212_sram_inv[0:1]),
		.out(chany_bottom_out[114]));

	mux_2level_tapbuf_size2 mux_bottom_track_231 (
		.in({chanx_right_in[33], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_213_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_213_sram_inv[0:1]),
		.out(chany_bottom_out[115]));

	mux_2level_tapbuf_size2 mux_bottom_track_233 (
		.in({chanx_right_in[32], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_214_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_214_sram_inv[0:1]),
		.out(chany_bottom_out[116]));

	mux_2level_tapbuf_size2 mux_bottom_track_235 (
		.in({chanx_right_in[31], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_215_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_215_sram_inv[0:1]),
		.out(chany_bottom_out[117]));

	mux_2level_tapbuf_size2 mux_bottom_track_241 (
		.in({chanx_right_in[28], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_216_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_216_sram_inv[0:1]),
		.out(chany_bottom_out[120]));

	mux_2level_tapbuf_size2 mux_bottom_track_243 (
		.in({chanx_right_in[27], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_217_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_217_sram_inv[0:1]),
		.out(chany_bottom_out[121]));

	mux_2level_tapbuf_size2 mux_bottom_track_245 (
		.in({chanx_right_in[26], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_218_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_218_sram_inv[0:1]),
		.out(chany_bottom_out[122]));

	mux_2level_tapbuf_size2 mux_bottom_track_247 (
		.in({chanx_right_in[25], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_219_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_219_sram_inv[0:1]),
		.out(chany_bottom_out[123]));

	mux_2level_tapbuf_size2 mux_bottom_track_249 (
		.in({chanx_right_in[24], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_220_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_220_sram_inv[0:1]),
		.out(chany_bottom_out[124]));

	mux_2level_tapbuf_size2 mux_bottom_track_251 (
		.in({chanx_right_in[23], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_221_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_221_sram_inv[0:1]),
		.out(chany_bottom_out[125]));

	mux_2level_tapbuf_size2 mux_bottom_track_253 (
		.in({chanx_right_in[22], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_222_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_222_sram_inv[0:1]),
		.out(chany_bottom_out[126]));

	mux_2level_tapbuf_size2 mux_bottom_track_255 (
		.in({chanx_right_in[21], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_223_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_223_sram_inv[0:1]),
		.out(chany_bottom_out[127]));

	mux_2level_tapbuf_size2 mux_bottom_track_261 (
		.in({chanx_right_in[18], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_224_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_224_sram_inv[0:1]),
		.out(chany_bottom_out[130]));

	mux_2level_tapbuf_size2 mux_bottom_track_263 (
		.in({chanx_right_in[17], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_225_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_225_sram_inv[0:1]),
		.out(chany_bottom_out[131]));

	mux_2level_tapbuf_size2 mux_bottom_track_265 (
		.in({chanx_right_in[16], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_226_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_226_sram_inv[0:1]),
		.out(chany_bottom_out[132]));

	mux_2level_tapbuf_size2 mux_bottom_track_267 (
		.in({chanx_right_in[15], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_227_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_227_sram_inv[0:1]),
		.out(chany_bottom_out[133]));

	mux_2level_tapbuf_size2 mux_bottom_track_269 (
		.in({chanx_right_in[14], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_228_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_228_sram_inv[0:1]),
		.out(chany_bottom_out[134]));

	mux_2level_tapbuf_size2 mux_bottom_track_271 (
		.in({chanx_right_in[13], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_229_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_229_sram_inv[0:1]),
		.out(chany_bottom_out[135]));

	mux_2level_tapbuf_size2 mux_bottom_track_273 (
		.in({chanx_right_in[12], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_230_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_230_sram_inv[0:1]),
		.out(chany_bottom_out[136]));

	mux_2level_tapbuf_size2 mux_bottom_track_275 (
		.in({chanx_right_in[11], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_231_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_231_sram_inv[0:1]),
		.out(chany_bottom_out[137]));

	mux_2level_tapbuf_size2 mux_bottom_track_281 (
		.in({chanx_right_in[8], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_232_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_232_sram_inv[0:1]),
		.out(chany_bottom_out[140]));

	mux_2level_tapbuf_size2 mux_bottom_track_283 (
		.in({chanx_right_in[7], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_233_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_233_sram_inv[0:1]),
		.out(chany_bottom_out[141]));

	mux_2level_tapbuf_size2 mux_bottom_track_285 (
		.in({chanx_right_in[6], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_234_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_234_sram_inv[0:1]),
		.out(chany_bottom_out[142]));

	mux_2level_tapbuf_size2 mux_bottom_track_287 (
		.in({chanx_right_in[5], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_235_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_235_sram_inv[0:1]),
		.out(chany_bottom_out[143]));

	mux_2level_tapbuf_size2 mux_bottom_track_289 (
		.in({chanx_right_in[4], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_236_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_236_sram_inv[0:1]),
		.out(chany_bottom_out[144]));

	mux_2level_tapbuf_size2 mux_bottom_track_291 (
		.in({chanx_right_in[3], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_237_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_237_sram_inv[0:1]),
		.out(chany_bottom_out[145]));

	mux_2level_tapbuf_size2 mux_bottom_track_293 (
		.in({chanx_right_in[2], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_238_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_238_sram_inv[0:1]),
		.out(chany_bottom_out[146]));

	mux_2level_tapbuf_size2 mux_bottom_track_295 (
		.in({chanx_right_in[1], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_239_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_239_sram_inv[0:1]),
		.out(chany_bottom_out[147]));

	mux_2level_tapbuf_size2_mem mem_right_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_0_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_1_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_2_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_6 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_3_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_4_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_5_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_6_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_14 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_7_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_8_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_22 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_9_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_10_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_11_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_12_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_30 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_13_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_14_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_34 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_15_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_16_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_17_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_18_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_46 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_19_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_20_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_21_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_52 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_22_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_54 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_23_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_24_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_62 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_25_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_26_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_27_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_28_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_70 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_29_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_30_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_31_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_32_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_33_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_34_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_86 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_35_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_36_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_37_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_38_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_94 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_39_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_40_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_102 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_41_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_42_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_106 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_43_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_44_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_110 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_45_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_46_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_47_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_48_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_49_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_124 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_50_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_126 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_51_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_52_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_53_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_54_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_134 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_55_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_56_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_142 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_57_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_58_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_59_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_60_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_60_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_150 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_61_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_61_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_62_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_62_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_63_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_63_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_64_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_64_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_65_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_65_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_66_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_66_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_166 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_67_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_67_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_68_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_68_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_69_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_69_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_70_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_70_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_174 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_71_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_71_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_72_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_72_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_182 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_73_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_73_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_74_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_74_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_75_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_75_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_76_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_76_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_190 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_77_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_77_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_78_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_78_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_78_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_79_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_79_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_79_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_79_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_80_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_80_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_80_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_80_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_81_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_81_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_81_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_81_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_82_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_82_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_82_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_206 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_82_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_83_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_83_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_83_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_83_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_84_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_84_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_84_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_210 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_84_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_85_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_85_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_85_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_212 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_85_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_86_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_86_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_86_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_214 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_86_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_87_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_87_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_87_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_220 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_87_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_88_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_88_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_88_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_222 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_88_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_89_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_89_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_89_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_89_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_90_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_90_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_90_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_226 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_90_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_91_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_91_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_91_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_228 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_91_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_92_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_92_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_92_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_230 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_92_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_93_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_93_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_93_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_93_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_94_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_94_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_94_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_234 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_94_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_95_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_95_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_95_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_95_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_96_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_96_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_96_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_242 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_96_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_97_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_97_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_97_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_244 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_97_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_98_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_98_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_98_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_246 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_98_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_99_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_99_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_99_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_99_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_100_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_100_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_100_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_250 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_100_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_101_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_101_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_101_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_252 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_101_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_102_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_102_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_102_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_254 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_102_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_103_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_103_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_103_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_260 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_103_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_104_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_104_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_104_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_262 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_104_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_105_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_105_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_105_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_105_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_106_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_106_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_106_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_266 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_106_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_107_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_107_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_107_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_268 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_107_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_108_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_108_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_108_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_270 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_108_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_109_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_109_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_109_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_109_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_110_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_110_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_110_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_274 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_110_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_111_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_111_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_111_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_111_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_112_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_112_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_112_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_282 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_112_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_113_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_113_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_113_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_284 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_113_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_114_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_114_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_114_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_286 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_114_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_115_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_115_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_115_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_115_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_116_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_116_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_116_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_290 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_116_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_117_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_117_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_117_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_292 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_117_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_118_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_118_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_118_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_294 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_118_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_119_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_119_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_119_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_119_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_120_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_120_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_120_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_3 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_120_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_121_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_121_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_121_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_5 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_121_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_122_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_122_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_122_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_7 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_122_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_123_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_123_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_123_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_123_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_124_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_124_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_124_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_11 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_124_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_125_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_125_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_125_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_13 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_125_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_126_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_126_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_126_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_15 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_126_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_127_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_127_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_127_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_21 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_127_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_128_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_128_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_128_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_23 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_128_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_129_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_129_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_129_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_129_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_130_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_130_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_130_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_27 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_130_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_131_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_131_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_131_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_29 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_131_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_132_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_132_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_132_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_31 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_132_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_133_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_133_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_133_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_133_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_134_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_134_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_134_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_35 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_134_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_135_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_135_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_135_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_135_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_136_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_136_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_136_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_43 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_136_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_137_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_137_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_137_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_45 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_137_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_138_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_138_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_138_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_47 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_138_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_139_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_139_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_139_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_139_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_140_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_140_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_140_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_51 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_140_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_141_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_141_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_141_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_53 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_141_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_142_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_142_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_142_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_55 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_142_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_143_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_143_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_143_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_61 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_143_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_144_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_144_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_144_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_63 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_144_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_145_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_145_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_145_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_145_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_146_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_146_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_146_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_67 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_146_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_147_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_147_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_147_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_69 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_147_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_148_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_148_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_148_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_71 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_148_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_149_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_149_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_149_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_149_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_150_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_150_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_150_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_75 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_150_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_151_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_151_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_151_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_151_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_152_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_152_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_152_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_83 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_152_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_153_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_153_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_153_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_85 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_153_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_154_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_154_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_154_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_87 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_154_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_155_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_155_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_155_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_155_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_156_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_156_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_156_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_91 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_156_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_157_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_157_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_157_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_93 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_157_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_158_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_158_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_158_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_95 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_158_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_159_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_159_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_159_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_101 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_159_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_160_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_160_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_160_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_103 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_160_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_161_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_161_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_161_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_105 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_161_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_162_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_162_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_162_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_107 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_162_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_163_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_163_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_163_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_109 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_163_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_164_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_164_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_164_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_111 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_164_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_165_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_165_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_165_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_113 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_165_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_166_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_166_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_166_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_115 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_166_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_167_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_167_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_167_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_121 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_167_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_168_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_168_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_168_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_123 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_168_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_169_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_169_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_169_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_125 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_169_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_170_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_170_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_170_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_127 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_170_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_171_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_171_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_171_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_129 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_171_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_172_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_172_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_172_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_131 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_172_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_173_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_173_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_173_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_133 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_173_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_174_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_174_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_174_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_135 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_174_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_175_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_175_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_175_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_141 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_175_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_176_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_176_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_176_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_143 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_176_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_177_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_177_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_177_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_145 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_177_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_178_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_178_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_178_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_147 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_178_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_179_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_179_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_179_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_149 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_179_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_180_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_180_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_180_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_151 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_180_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_181_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_181_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_181_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_153 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_181_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_182_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_182_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_182_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_155 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_182_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_183_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_183_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_183_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_161 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_183_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_184_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_184_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_184_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_163 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_184_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_185_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_185_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_185_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_165 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_185_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_186_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_186_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_186_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_167 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_186_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_187_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_187_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_187_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_169 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_187_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_188_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_188_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_188_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_171 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_188_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_189_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_189_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_189_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_173 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_189_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_190_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_190_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_190_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_175 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_190_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_191_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_191_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_191_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_181 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_191_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_192_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_192_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_192_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_183 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_192_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_193_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_193_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_193_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_185 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_193_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_194_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_194_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_194_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_187 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_194_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_195_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_195_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_195_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_189 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_195_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_196_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_196_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_196_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_191 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_196_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_197_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_197_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_197_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_193 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_197_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_198_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_198_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_198_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_195 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_198_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_199_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_199_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_199_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_201 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_199_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_200_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_200_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_200_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_203 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_200_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_201_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_201_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_201_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_205 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_201_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_202_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_202_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_202_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_207 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_202_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_203_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_203_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_203_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_209 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_203_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_204_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_204_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_204_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_211 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_204_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_205_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_205_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_205_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_213 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_205_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_206_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_206_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_206_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_215 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_206_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_207_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_207_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_207_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_221 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_207_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_208_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_208_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_208_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_223 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_208_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_209_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_209_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_209_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_225 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_209_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_210_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_210_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_210_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_227 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_210_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_211_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_211_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_211_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_229 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_211_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_212_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_212_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_212_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_231 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_212_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_213_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_213_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_213_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_233 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_213_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_214_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_214_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_214_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_235 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_214_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_215_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_215_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_215_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_241 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_215_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_216_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_216_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_216_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_243 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_216_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_217_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_217_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_217_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_245 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_217_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_218_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_218_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_218_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_247 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_218_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_219_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_219_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_219_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_249 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_219_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_220_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_220_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_220_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_251 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_220_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_221_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_221_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_221_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_253 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_221_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_222_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_222_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_222_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_255 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_222_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_223_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_223_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_223_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_261 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_223_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_224_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_224_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_224_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_263 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_224_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_225_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_225_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_225_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_265 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_225_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_226_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_226_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_226_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_267 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_226_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_227_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_227_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_227_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_269 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_227_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_228_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_228_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_228_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_271 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_228_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_229_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_229_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_229_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_273 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_229_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_230_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_230_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_230_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_275 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_230_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_231_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_231_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_231_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_281 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_231_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_232_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_232_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_232_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_283 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_232_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_233_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_233_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_233_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_285 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_233_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_234_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_234_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_234_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_287 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_234_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_235_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_235_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_235_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_289 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_235_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_236_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_236_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_236_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_291 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_236_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_237_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_237_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_237_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_293 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_237_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_238_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_238_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_238_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_295 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_238_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_239_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_239_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_0__11_ -----

//----- Default net type -----
`default_nettype wire



