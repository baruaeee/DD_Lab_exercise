//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[11][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Mon Jul  7 22:55:54 2025
//-------------------------------------------
//----- Default net type -----
// `default_nettype none

// ----- Verilog module for sb_11__0_ -----
module sb_11__0_(pReset,
                 prog_clk,
                 chany_top_in,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_,
                 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
                 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                 chanx_left_in,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_,
                 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                 ccff_head,
                 chany_top_out,
                 chanx_left_out,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:149] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:149] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:149] chany_top_out;
//----- OUTPUT PORTS -----
output [0:149] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_2level_tapbuf_size2_0_sram;
wire [0:1] mux_2level_tapbuf_size2_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_10_sram;
wire [0:1] mux_2level_tapbuf_size2_10_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_11_sram;
wire [0:1] mux_2level_tapbuf_size2_11_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_12_sram;
wire [0:1] mux_2level_tapbuf_size2_12_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_13_sram;
wire [0:1] mux_2level_tapbuf_size2_13_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_14_sram;
wire [0:1] mux_2level_tapbuf_size2_14_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_15_sram;
wire [0:1] mux_2level_tapbuf_size2_15_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_16_sram;
wire [0:1] mux_2level_tapbuf_size2_16_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_17_sram;
wire [0:1] mux_2level_tapbuf_size2_17_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_18_sram;
wire [0:1] mux_2level_tapbuf_size2_18_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_19_sram;
wire [0:1] mux_2level_tapbuf_size2_19_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_1_sram;
wire [0:1] mux_2level_tapbuf_size2_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_20_sram;
wire [0:1] mux_2level_tapbuf_size2_20_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_21_sram;
wire [0:1] mux_2level_tapbuf_size2_21_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_22_sram;
wire [0:1] mux_2level_tapbuf_size2_22_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_23_sram;
wire [0:1] mux_2level_tapbuf_size2_23_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_24_sram;
wire [0:1] mux_2level_tapbuf_size2_24_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_25_sram;
wire [0:1] mux_2level_tapbuf_size2_25_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_26_sram;
wire [0:1] mux_2level_tapbuf_size2_26_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_27_sram;
wire [0:1] mux_2level_tapbuf_size2_27_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_28_sram;
wire [0:1] mux_2level_tapbuf_size2_28_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_29_sram;
wire [0:1] mux_2level_tapbuf_size2_29_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_2_sram;
wire [0:1] mux_2level_tapbuf_size2_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_30_sram;
wire [0:1] mux_2level_tapbuf_size2_30_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_31_sram;
wire [0:1] mux_2level_tapbuf_size2_31_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_32_sram;
wire [0:1] mux_2level_tapbuf_size2_32_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_33_sram;
wire [0:1] mux_2level_tapbuf_size2_33_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_34_sram;
wire [0:1] mux_2level_tapbuf_size2_34_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_35_sram;
wire [0:1] mux_2level_tapbuf_size2_35_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_36_sram;
wire [0:1] mux_2level_tapbuf_size2_36_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_37_sram;
wire [0:1] mux_2level_tapbuf_size2_37_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_38_sram;
wire [0:1] mux_2level_tapbuf_size2_38_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_39_sram;
wire [0:1] mux_2level_tapbuf_size2_39_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_3_sram;
wire [0:1] mux_2level_tapbuf_size2_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_40_sram;
wire [0:1] mux_2level_tapbuf_size2_40_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_41_sram;
wire [0:1] mux_2level_tapbuf_size2_41_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_42_sram;
wire [0:1] mux_2level_tapbuf_size2_42_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_43_sram;
wire [0:1] mux_2level_tapbuf_size2_43_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_44_sram;
wire [0:1] mux_2level_tapbuf_size2_44_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_45_sram;
wire [0:1] mux_2level_tapbuf_size2_45_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_46_sram;
wire [0:1] mux_2level_tapbuf_size2_46_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_47_sram;
wire [0:1] mux_2level_tapbuf_size2_47_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_48_sram;
wire [0:1] mux_2level_tapbuf_size2_48_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_49_sram;
wire [0:1] mux_2level_tapbuf_size2_49_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_4_sram;
wire [0:1] mux_2level_tapbuf_size2_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_50_sram;
wire [0:1] mux_2level_tapbuf_size2_50_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_51_sram;
wire [0:1] mux_2level_tapbuf_size2_51_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_52_sram;
wire [0:1] mux_2level_tapbuf_size2_52_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_53_sram;
wire [0:1] mux_2level_tapbuf_size2_53_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_54_sram;
wire [0:1] mux_2level_tapbuf_size2_54_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_55_sram;
wire [0:1] mux_2level_tapbuf_size2_55_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_56_sram;
wire [0:1] mux_2level_tapbuf_size2_56_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_57_sram;
wire [0:1] mux_2level_tapbuf_size2_57_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_58_sram;
wire [0:1] mux_2level_tapbuf_size2_58_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_59_sram;
wire [0:1] mux_2level_tapbuf_size2_59_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_5_sram;
wire [0:1] mux_2level_tapbuf_size2_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_6_sram;
wire [0:1] mux_2level_tapbuf_size2_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_7_sram;
wire [0:1] mux_2level_tapbuf_size2_7_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_8_sram;
wire [0:1] mux_2level_tapbuf_size2_8_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_9_sram;
wire [0:1] mux_2level_tapbuf_size2_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_9_ccff_tail;
wire [0:1] mux_2level_tapbuf_size3_0_sram;
wire [0:1] mux_2level_tapbuf_size3_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_100_sram;
wire [0:1] mux_2level_tapbuf_size3_100_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_101_sram;
wire [0:1] mux_2level_tapbuf_size3_101_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_102_sram;
wire [0:1] mux_2level_tapbuf_size3_102_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_103_sram;
wire [0:1] mux_2level_tapbuf_size3_103_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_104_sram;
wire [0:1] mux_2level_tapbuf_size3_104_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_105_sram;
wire [0:1] mux_2level_tapbuf_size3_105_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_106_sram;
wire [0:1] mux_2level_tapbuf_size3_106_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_107_sram;
wire [0:1] mux_2level_tapbuf_size3_107_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_108_sram;
wire [0:1] mux_2level_tapbuf_size3_108_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_109_sram;
wire [0:1] mux_2level_tapbuf_size3_109_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_10_sram;
wire [0:1] mux_2level_tapbuf_size3_10_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_110_sram;
wire [0:1] mux_2level_tapbuf_size3_110_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_111_sram;
wire [0:1] mux_2level_tapbuf_size3_111_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_112_sram;
wire [0:1] mux_2level_tapbuf_size3_112_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_113_sram;
wire [0:1] mux_2level_tapbuf_size3_113_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_114_sram;
wire [0:1] mux_2level_tapbuf_size3_114_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_115_sram;
wire [0:1] mux_2level_tapbuf_size3_115_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_116_sram;
wire [0:1] mux_2level_tapbuf_size3_116_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_117_sram;
wire [0:1] mux_2level_tapbuf_size3_117_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_118_sram;
wire [0:1] mux_2level_tapbuf_size3_118_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_119_sram;
wire [0:1] mux_2level_tapbuf_size3_119_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_11_sram;
wire [0:1] mux_2level_tapbuf_size3_11_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_120_sram;
wire [0:1] mux_2level_tapbuf_size3_120_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_121_sram;
wire [0:1] mux_2level_tapbuf_size3_121_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_122_sram;
wire [0:1] mux_2level_tapbuf_size3_122_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_123_sram;
wire [0:1] mux_2level_tapbuf_size3_123_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_124_sram;
wire [0:1] mux_2level_tapbuf_size3_124_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_125_sram;
wire [0:1] mux_2level_tapbuf_size3_125_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_126_sram;
wire [0:1] mux_2level_tapbuf_size3_126_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_127_sram;
wire [0:1] mux_2level_tapbuf_size3_127_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_128_sram;
wire [0:1] mux_2level_tapbuf_size3_128_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_129_sram;
wire [0:1] mux_2level_tapbuf_size3_129_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_12_sram;
wire [0:1] mux_2level_tapbuf_size3_12_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_130_sram;
wire [0:1] mux_2level_tapbuf_size3_130_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_131_sram;
wire [0:1] mux_2level_tapbuf_size3_131_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_132_sram;
wire [0:1] mux_2level_tapbuf_size3_132_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_133_sram;
wire [0:1] mux_2level_tapbuf_size3_133_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_134_sram;
wire [0:1] mux_2level_tapbuf_size3_134_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_135_sram;
wire [0:1] mux_2level_tapbuf_size3_135_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_136_sram;
wire [0:1] mux_2level_tapbuf_size3_136_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_137_sram;
wire [0:1] mux_2level_tapbuf_size3_137_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_138_sram;
wire [0:1] mux_2level_tapbuf_size3_138_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_139_sram;
wire [0:1] mux_2level_tapbuf_size3_139_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_13_sram;
wire [0:1] mux_2level_tapbuf_size3_13_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_140_sram;
wire [0:1] mux_2level_tapbuf_size3_140_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_141_sram;
wire [0:1] mux_2level_tapbuf_size3_141_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_142_sram;
wire [0:1] mux_2level_tapbuf_size3_142_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_143_sram;
wire [0:1] mux_2level_tapbuf_size3_143_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_144_sram;
wire [0:1] mux_2level_tapbuf_size3_144_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_145_sram;
wire [0:1] mux_2level_tapbuf_size3_145_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_146_sram;
wire [0:1] mux_2level_tapbuf_size3_146_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_147_sram;
wire [0:1] mux_2level_tapbuf_size3_147_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_148_sram;
wire [0:1] mux_2level_tapbuf_size3_148_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_149_sram;
wire [0:1] mux_2level_tapbuf_size3_149_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_14_sram;
wire [0:1] mux_2level_tapbuf_size3_14_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_150_sram;
wire [0:1] mux_2level_tapbuf_size3_150_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_151_sram;
wire [0:1] mux_2level_tapbuf_size3_151_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_152_sram;
wire [0:1] mux_2level_tapbuf_size3_152_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_153_sram;
wire [0:1] mux_2level_tapbuf_size3_153_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_154_sram;
wire [0:1] mux_2level_tapbuf_size3_154_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_155_sram;
wire [0:1] mux_2level_tapbuf_size3_155_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_156_sram;
wire [0:1] mux_2level_tapbuf_size3_156_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_157_sram;
wire [0:1] mux_2level_tapbuf_size3_157_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_158_sram;
wire [0:1] mux_2level_tapbuf_size3_158_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_159_sram;
wire [0:1] mux_2level_tapbuf_size3_159_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_15_sram;
wire [0:1] mux_2level_tapbuf_size3_15_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_160_sram;
wire [0:1] mux_2level_tapbuf_size3_160_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_161_sram;
wire [0:1] mux_2level_tapbuf_size3_161_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_162_sram;
wire [0:1] mux_2level_tapbuf_size3_162_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_163_sram;
wire [0:1] mux_2level_tapbuf_size3_163_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_164_sram;
wire [0:1] mux_2level_tapbuf_size3_164_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_165_sram;
wire [0:1] mux_2level_tapbuf_size3_165_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_166_sram;
wire [0:1] mux_2level_tapbuf_size3_166_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_167_sram;
wire [0:1] mux_2level_tapbuf_size3_167_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_168_sram;
wire [0:1] mux_2level_tapbuf_size3_168_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_169_sram;
wire [0:1] mux_2level_tapbuf_size3_169_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_16_sram;
wire [0:1] mux_2level_tapbuf_size3_16_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_170_sram;
wire [0:1] mux_2level_tapbuf_size3_170_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_171_sram;
wire [0:1] mux_2level_tapbuf_size3_171_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_172_sram;
wire [0:1] mux_2level_tapbuf_size3_172_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_173_sram;
wire [0:1] mux_2level_tapbuf_size3_173_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_174_sram;
wire [0:1] mux_2level_tapbuf_size3_174_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_175_sram;
wire [0:1] mux_2level_tapbuf_size3_175_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_176_sram;
wire [0:1] mux_2level_tapbuf_size3_176_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_177_sram;
wire [0:1] mux_2level_tapbuf_size3_177_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_178_sram;
wire [0:1] mux_2level_tapbuf_size3_178_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_179_sram;
wire [0:1] mux_2level_tapbuf_size3_179_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_17_sram;
wire [0:1] mux_2level_tapbuf_size3_17_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_180_sram;
wire [0:1] mux_2level_tapbuf_size3_180_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_181_sram;
wire [0:1] mux_2level_tapbuf_size3_181_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_182_sram;
wire [0:1] mux_2level_tapbuf_size3_182_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_183_sram;
wire [0:1] mux_2level_tapbuf_size3_183_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_184_sram;
wire [0:1] mux_2level_tapbuf_size3_184_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_185_sram;
wire [0:1] mux_2level_tapbuf_size3_185_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_186_sram;
wire [0:1] mux_2level_tapbuf_size3_186_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_187_sram;
wire [0:1] mux_2level_tapbuf_size3_187_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_188_sram;
wire [0:1] mux_2level_tapbuf_size3_188_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_189_sram;
wire [0:1] mux_2level_tapbuf_size3_189_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_18_sram;
wire [0:1] mux_2level_tapbuf_size3_18_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_190_sram;
wire [0:1] mux_2level_tapbuf_size3_190_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_191_sram;
wire [0:1] mux_2level_tapbuf_size3_191_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_192_sram;
wire [0:1] mux_2level_tapbuf_size3_192_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_193_sram;
wire [0:1] mux_2level_tapbuf_size3_193_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_194_sram;
wire [0:1] mux_2level_tapbuf_size3_194_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_195_sram;
wire [0:1] mux_2level_tapbuf_size3_195_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_196_sram;
wire [0:1] mux_2level_tapbuf_size3_196_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_197_sram;
wire [0:1] mux_2level_tapbuf_size3_197_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_198_sram;
wire [0:1] mux_2level_tapbuf_size3_198_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_199_sram;
wire [0:1] mux_2level_tapbuf_size3_199_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_19_sram;
wire [0:1] mux_2level_tapbuf_size3_19_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_1_sram;
wire [0:1] mux_2level_tapbuf_size3_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_200_sram;
wire [0:1] mux_2level_tapbuf_size3_200_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_201_sram;
wire [0:1] mux_2level_tapbuf_size3_201_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_202_sram;
wire [0:1] mux_2level_tapbuf_size3_202_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_203_sram;
wire [0:1] mux_2level_tapbuf_size3_203_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_204_sram;
wire [0:1] mux_2level_tapbuf_size3_204_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_205_sram;
wire [0:1] mux_2level_tapbuf_size3_205_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_206_sram;
wire [0:1] mux_2level_tapbuf_size3_206_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_207_sram;
wire [0:1] mux_2level_tapbuf_size3_207_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_208_sram;
wire [0:1] mux_2level_tapbuf_size3_208_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_209_sram;
wire [0:1] mux_2level_tapbuf_size3_209_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_20_sram;
wire [0:1] mux_2level_tapbuf_size3_20_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_210_sram;
wire [0:1] mux_2level_tapbuf_size3_210_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_211_sram;
wire [0:1] mux_2level_tapbuf_size3_211_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_212_sram;
wire [0:1] mux_2level_tapbuf_size3_212_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_213_sram;
wire [0:1] mux_2level_tapbuf_size3_213_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_214_sram;
wire [0:1] mux_2level_tapbuf_size3_214_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_215_sram;
wire [0:1] mux_2level_tapbuf_size3_215_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_216_sram;
wire [0:1] mux_2level_tapbuf_size3_216_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_217_sram;
wire [0:1] mux_2level_tapbuf_size3_217_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_218_sram;
wire [0:1] mux_2level_tapbuf_size3_218_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_219_sram;
wire [0:1] mux_2level_tapbuf_size3_219_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_21_sram;
wire [0:1] mux_2level_tapbuf_size3_21_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_220_sram;
wire [0:1] mux_2level_tapbuf_size3_220_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_221_sram;
wire [0:1] mux_2level_tapbuf_size3_221_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_222_sram;
wire [0:1] mux_2level_tapbuf_size3_222_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_223_sram;
wire [0:1] mux_2level_tapbuf_size3_223_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_224_sram;
wire [0:1] mux_2level_tapbuf_size3_224_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_225_sram;
wire [0:1] mux_2level_tapbuf_size3_225_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_226_sram;
wire [0:1] mux_2level_tapbuf_size3_226_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_227_sram;
wire [0:1] mux_2level_tapbuf_size3_227_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_228_sram;
wire [0:1] mux_2level_tapbuf_size3_228_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_229_sram;
wire [0:1] mux_2level_tapbuf_size3_229_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_22_sram;
wire [0:1] mux_2level_tapbuf_size3_22_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_230_sram;
wire [0:1] mux_2level_tapbuf_size3_230_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_231_sram;
wire [0:1] mux_2level_tapbuf_size3_231_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_232_sram;
wire [0:1] mux_2level_tapbuf_size3_232_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_233_sram;
wire [0:1] mux_2level_tapbuf_size3_233_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_234_sram;
wire [0:1] mux_2level_tapbuf_size3_234_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_235_sram;
wire [0:1] mux_2level_tapbuf_size3_235_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_236_sram;
wire [0:1] mux_2level_tapbuf_size3_236_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_237_sram;
wire [0:1] mux_2level_tapbuf_size3_237_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_238_sram;
wire [0:1] mux_2level_tapbuf_size3_238_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_239_sram;
wire [0:1] mux_2level_tapbuf_size3_239_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_23_sram;
wire [0:1] mux_2level_tapbuf_size3_23_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_24_sram;
wire [0:1] mux_2level_tapbuf_size3_24_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_25_sram;
wire [0:1] mux_2level_tapbuf_size3_25_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_26_sram;
wire [0:1] mux_2level_tapbuf_size3_26_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_27_sram;
wire [0:1] mux_2level_tapbuf_size3_27_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_28_sram;
wire [0:1] mux_2level_tapbuf_size3_28_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_29_sram;
wire [0:1] mux_2level_tapbuf_size3_29_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_2_sram;
wire [0:1] mux_2level_tapbuf_size3_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_30_sram;
wire [0:1] mux_2level_tapbuf_size3_30_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_31_sram;
wire [0:1] mux_2level_tapbuf_size3_31_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_32_sram;
wire [0:1] mux_2level_tapbuf_size3_32_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_33_sram;
wire [0:1] mux_2level_tapbuf_size3_33_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_34_sram;
wire [0:1] mux_2level_tapbuf_size3_34_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_35_sram;
wire [0:1] mux_2level_tapbuf_size3_35_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_36_sram;
wire [0:1] mux_2level_tapbuf_size3_36_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_37_sram;
wire [0:1] mux_2level_tapbuf_size3_37_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_38_sram;
wire [0:1] mux_2level_tapbuf_size3_38_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_39_sram;
wire [0:1] mux_2level_tapbuf_size3_39_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_3_sram;
wire [0:1] mux_2level_tapbuf_size3_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_40_sram;
wire [0:1] mux_2level_tapbuf_size3_40_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_41_sram;
wire [0:1] mux_2level_tapbuf_size3_41_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_42_sram;
wire [0:1] mux_2level_tapbuf_size3_42_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_43_sram;
wire [0:1] mux_2level_tapbuf_size3_43_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_44_sram;
wire [0:1] mux_2level_tapbuf_size3_44_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_45_sram;
wire [0:1] mux_2level_tapbuf_size3_45_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_46_sram;
wire [0:1] mux_2level_tapbuf_size3_46_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_47_sram;
wire [0:1] mux_2level_tapbuf_size3_47_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_48_sram;
wire [0:1] mux_2level_tapbuf_size3_48_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_49_sram;
wire [0:1] mux_2level_tapbuf_size3_49_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_4_sram;
wire [0:1] mux_2level_tapbuf_size3_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_50_sram;
wire [0:1] mux_2level_tapbuf_size3_50_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_51_sram;
wire [0:1] mux_2level_tapbuf_size3_51_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_52_sram;
wire [0:1] mux_2level_tapbuf_size3_52_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_53_sram;
wire [0:1] mux_2level_tapbuf_size3_53_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_54_sram;
wire [0:1] mux_2level_tapbuf_size3_54_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_55_sram;
wire [0:1] mux_2level_tapbuf_size3_55_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_56_sram;
wire [0:1] mux_2level_tapbuf_size3_56_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_57_sram;
wire [0:1] mux_2level_tapbuf_size3_57_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_58_sram;
wire [0:1] mux_2level_tapbuf_size3_58_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_59_sram;
wire [0:1] mux_2level_tapbuf_size3_59_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_5_sram;
wire [0:1] mux_2level_tapbuf_size3_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_60_sram;
wire [0:1] mux_2level_tapbuf_size3_60_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_61_sram;
wire [0:1] mux_2level_tapbuf_size3_61_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_62_sram;
wire [0:1] mux_2level_tapbuf_size3_62_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_63_sram;
wire [0:1] mux_2level_tapbuf_size3_63_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_64_sram;
wire [0:1] mux_2level_tapbuf_size3_64_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_65_sram;
wire [0:1] mux_2level_tapbuf_size3_65_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_66_sram;
wire [0:1] mux_2level_tapbuf_size3_66_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_67_sram;
wire [0:1] mux_2level_tapbuf_size3_67_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_68_sram;
wire [0:1] mux_2level_tapbuf_size3_68_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_69_sram;
wire [0:1] mux_2level_tapbuf_size3_69_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_6_sram;
wire [0:1] mux_2level_tapbuf_size3_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_70_sram;
wire [0:1] mux_2level_tapbuf_size3_70_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_71_sram;
wire [0:1] mux_2level_tapbuf_size3_71_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_72_sram;
wire [0:1] mux_2level_tapbuf_size3_72_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_73_sram;
wire [0:1] mux_2level_tapbuf_size3_73_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_74_sram;
wire [0:1] mux_2level_tapbuf_size3_74_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_75_sram;
wire [0:1] mux_2level_tapbuf_size3_75_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_76_sram;
wire [0:1] mux_2level_tapbuf_size3_76_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_77_sram;
wire [0:1] mux_2level_tapbuf_size3_77_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_78_sram;
wire [0:1] mux_2level_tapbuf_size3_78_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_79_sram;
wire [0:1] mux_2level_tapbuf_size3_79_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_7_sram;
wire [0:1] mux_2level_tapbuf_size3_7_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_80_sram;
wire [0:1] mux_2level_tapbuf_size3_80_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_81_sram;
wire [0:1] mux_2level_tapbuf_size3_81_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_82_sram;
wire [0:1] mux_2level_tapbuf_size3_82_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_83_sram;
wire [0:1] mux_2level_tapbuf_size3_83_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_84_sram;
wire [0:1] mux_2level_tapbuf_size3_84_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_85_sram;
wire [0:1] mux_2level_tapbuf_size3_85_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_86_sram;
wire [0:1] mux_2level_tapbuf_size3_86_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_87_sram;
wire [0:1] mux_2level_tapbuf_size3_87_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_88_sram;
wire [0:1] mux_2level_tapbuf_size3_88_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_89_sram;
wire [0:1] mux_2level_tapbuf_size3_89_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_8_sram;
wire [0:1] mux_2level_tapbuf_size3_8_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_90_sram;
wire [0:1] mux_2level_tapbuf_size3_90_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_91_sram;
wire [0:1] mux_2level_tapbuf_size3_91_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_92_sram;
wire [0:1] mux_2level_tapbuf_size3_92_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_93_sram;
wire [0:1] mux_2level_tapbuf_size3_93_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_94_sram;
wire [0:1] mux_2level_tapbuf_size3_94_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_95_sram;
wire [0:1] mux_2level_tapbuf_size3_95_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_96_sram;
wire [0:1] mux_2level_tapbuf_size3_96_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_97_sram;
wire [0:1] mux_2level_tapbuf_size3_97_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_98_sram;
wire [0:1] mux_2level_tapbuf_size3_98_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_99_sram;
wire [0:1] mux_2level_tapbuf_size3_99_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_9_sram;
wire [0:1] mux_2level_tapbuf_size3_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_100_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_101_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_102_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_103_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_104_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_105_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_106_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_107_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_108_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_109_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_110_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_111_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_112_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_113_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_114_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_115_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_116_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_117_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_118_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_119_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_120_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_121_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_122_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_123_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_124_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_125_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_126_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_127_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_128_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_129_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_130_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_131_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_132_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_133_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_134_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_135_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_136_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_137_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_138_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_139_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_140_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_141_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_142_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_143_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_144_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_145_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_146_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_147_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_148_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_149_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_150_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_151_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_152_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_153_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_154_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_155_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_156_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_157_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_158_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_159_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_160_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_161_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_162_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_163_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_164_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_165_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_166_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_167_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_168_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_169_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_170_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_171_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_172_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_173_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_174_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_175_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_176_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_177_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_178_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_179_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_180_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_181_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_182_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_183_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_184_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_185_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_186_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_187_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_188_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_189_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_190_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_191_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_192_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_193_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_194_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_195_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_196_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_197_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_198_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_199_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_200_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_201_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_202_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_203_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_204_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_205_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_206_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_207_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_208_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_209_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_210_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_211_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_212_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_213_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_214_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_215_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_216_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_217_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_218_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_219_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_220_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_221_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_222_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_223_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_224_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_225_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_226_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_227_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_228_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_229_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_230_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_231_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_232_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_233_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_234_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_235_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_236_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_237_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_238_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_239_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_79_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_80_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_81_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_82_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_83_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_84_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_85_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_86_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_87_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_88_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_89_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_90_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_91_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_92_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_93_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_94_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_95_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_96_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_97_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_98_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_99_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size3 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[0]}),
		.sram(mux_2level_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_0_sram_inv[0:1]),
		.out(chany_top_out[0]));

	mux_2level_tapbuf_size3 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[149]}),
		.sram(mux_2level_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_1_sram_inv[0:1]),
		.out(chany_top_out[1]));

	mux_2level_tapbuf_size3 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[148]}),
		.sram(mux_2level_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_2_sram_inv[0:1]),
		.out(chany_top_out[2]));

	mux_2level_tapbuf_size3 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[147]}),
		.sram(mux_2level_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_3_sram_inv[0:1]),
		.out(chany_top_out[3]));

	mux_2level_tapbuf_size3 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[146]}),
		.sram(mux_2level_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_4_sram_inv[0:1]),
		.out(chany_top_out[4]));

	mux_2level_tapbuf_size3 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[145]}),
		.sram(mux_2level_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_5_sram_inv[0:1]),
		.out(chany_top_out[5]));

	mux_2level_tapbuf_size3 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[144]}),
		.sram(mux_2level_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_6_sram_inv[0:1]),
		.out(chany_top_out[6]));

	mux_2level_tapbuf_size3 mux_top_track_14 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[143]}),
		.sram(mux_2level_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_7_sram_inv[0:1]),
		.out(chany_top_out[7]));

	mux_2level_tapbuf_size3 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[140]}),
		.sram(mux_2level_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_8_sram_inv[0:1]),
		.out(chany_top_out[10]));

	mux_2level_tapbuf_size3 mux_top_track_22 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[139]}),
		.sram(mux_2level_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_9_sram_inv[0:1]),
		.out(chany_top_out[11]));

	mux_2level_tapbuf_size3 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[138]}),
		.sram(mux_2level_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_10_sram_inv[0:1]),
		.out(chany_top_out[12]));

	mux_2level_tapbuf_size3 mux_top_track_26 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[137]}),
		.sram(mux_2level_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_11_sram_inv[0:1]),
		.out(chany_top_out[13]));

	mux_2level_tapbuf_size3 mux_top_track_28 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[136]}),
		.sram(mux_2level_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_12_sram_inv[0:1]),
		.out(chany_top_out[14]));

	mux_2level_tapbuf_size3 mux_top_track_30 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[135]}),
		.sram(mux_2level_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_13_sram_inv[0:1]),
		.out(chany_top_out[15]));

	mux_2level_tapbuf_size3 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[134]}),
		.sram(mux_2level_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_14_sram_inv[0:1]),
		.out(chany_top_out[16]));

	mux_2level_tapbuf_size3 mux_top_track_34 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[133]}),
		.sram(mux_2level_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_15_sram_inv[0:1]),
		.out(chany_top_out[17]));

	mux_2level_tapbuf_size3 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[130]}),
		.sram(mux_2level_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_16_sram_inv[0:1]),
		.out(chany_top_out[20]));

	mux_2level_tapbuf_size3 mux_top_track_42 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[129]}),
		.sram(mux_2level_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_17_sram_inv[0:1]),
		.out(chany_top_out[21]));

	mux_2level_tapbuf_size3 mux_top_track_44 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[128]}),
		.sram(mux_2level_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_18_sram_inv[0:1]),
		.out(chany_top_out[22]));

	mux_2level_tapbuf_size3 mux_top_track_46 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[127]}),
		.sram(mux_2level_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_19_sram_inv[0:1]),
		.out(chany_top_out[23]));

	mux_2level_tapbuf_size3 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[126]}),
		.sram(mux_2level_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_20_sram_inv[0:1]),
		.out(chany_top_out[24]));

	mux_2level_tapbuf_size3 mux_top_track_50 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[125]}),
		.sram(mux_2level_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_21_sram_inv[0:1]),
		.out(chany_top_out[25]));

	mux_2level_tapbuf_size3 mux_top_track_52 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[124]}),
		.sram(mux_2level_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_22_sram_inv[0:1]),
		.out(chany_top_out[26]));

	mux_2level_tapbuf_size3 mux_top_track_54 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[123]}),
		.sram(mux_2level_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_23_sram_inv[0:1]),
		.out(chany_top_out[27]));

	mux_2level_tapbuf_size3 mux_top_track_60 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[120]}),
		.sram(mux_2level_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_24_sram_inv[0:1]),
		.out(chany_top_out[30]));

	mux_2level_tapbuf_size3 mux_top_track_62 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[119]}),
		.sram(mux_2level_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_25_sram_inv[0:1]),
		.out(chany_top_out[31]));

	mux_2level_tapbuf_size3 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[118]}),
		.sram(mux_2level_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_26_sram_inv[0:1]),
		.out(chany_top_out[32]));

	mux_2level_tapbuf_size3 mux_top_track_66 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[117]}),
		.sram(mux_2level_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_27_sram_inv[0:1]),
		.out(chany_top_out[33]));

	mux_2level_tapbuf_size3 mux_top_track_68 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[116]}),
		.sram(mux_2level_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_28_sram_inv[0:1]),
		.out(chany_top_out[34]));

	mux_2level_tapbuf_size3 mux_top_track_70 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[115]}),
		.sram(mux_2level_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_29_sram_inv[0:1]),
		.out(chany_top_out[35]));

	mux_2level_tapbuf_size3 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[114]}),
		.sram(mux_2level_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_30_sram_inv[0:1]),
		.out(chany_top_out[36]));

	mux_2level_tapbuf_size3 mux_top_track_74 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[113]}),
		.sram(mux_2level_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_31_sram_inv[0:1]),
		.out(chany_top_out[37]));

	mux_2level_tapbuf_size3 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[110]}),
		.sram(mux_2level_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_32_sram_inv[0:1]),
		.out(chany_top_out[40]));

	mux_2level_tapbuf_size3 mux_top_track_82 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[109]}),
		.sram(mux_2level_tapbuf_size3_33_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_33_sram_inv[0:1]),
		.out(chany_top_out[41]));

	mux_2level_tapbuf_size3 mux_top_track_84 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[108]}),
		.sram(mux_2level_tapbuf_size3_34_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_34_sram_inv[0:1]),
		.out(chany_top_out[42]));

	mux_2level_tapbuf_size3 mux_top_track_86 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[107]}),
		.sram(mux_2level_tapbuf_size3_35_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_35_sram_inv[0:1]),
		.out(chany_top_out[43]));

	mux_2level_tapbuf_size3 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[106]}),
		.sram(mux_2level_tapbuf_size3_36_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_36_sram_inv[0:1]),
		.out(chany_top_out[44]));

	mux_2level_tapbuf_size3 mux_top_track_90 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[105]}),
		.sram(mux_2level_tapbuf_size3_37_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_37_sram_inv[0:1]),
		.out(chany_top_out[45]));

	mux_2level_tapbuf_size3 mux_top_track_92 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[104]}),
		.sram(mux_2level_tapbuf_size3_38_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_38_sram_inv[0:1]),
		.out(chany_top_out[46]));

	mux_2level_tapbuf_size3 mux_top_track_94 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[103]}),
		.sram(mux_2level_tapbuf_size3_39_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_39_sram_inv[0:1]),
		.out(chany_top_out[47]));

	mux_2level_tapbuf_size3 mux_top_track_100 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[100]}),
		.sram(mux_2level_tapbuf_size3_40_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_40_sram_inv[0:1]),
		.out(chany_top_out[50]));

	mux_2level_tapbuf_size3 mux_top_track_102 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[99]}),
		.sram(mux_2level_tapbuf_size3_41_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_41_sram_inv[0:1]),
		.out(chany_top_out[51]));

	mux_2level_tapbuf_size3 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[98]}),
		.sram(mux_2level_tapbuf_size3_42_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_42_sram_inv[0:1]),
		.out(chany_top_out[52]));

	mux_2level_tapbuf_size3 mux_top_track_106 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[97]}),
		.sram(mux_2level_tapbuf_size3_43_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_43_sram_inv[0:1]),
		.out(chany_top_out[53]));

	mux_2level_tapbuf_size3 mux_top_track_108 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[96]}),
		.sram(mux_2level_tapbuf_size3_44_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_44_sram_inv[0:1]),
		.out(chany_top_out[54]));

	mux_2level_tapbuf_size3 mux_top_track_110 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[95]}),
		.sram(mux_2level_tapbuf_size3_45_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_45_sram_inv[0:1]),
		.out(chany_top_out[55]));

	mux_2level_tapbuf_size3 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[94]}),
		.sram(mux_2level_tapbuf_size3_46_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_46_sram_inv[0:1]),
		.out(chany_top_out[56]));

	mux_2level_tapbuf_size3 mux_top_track_114 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[93]}),
		.sram(mux_2level_tapbuf_size3_47_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_47_sram_inv[0:1]),
		.out(chany_top_out[57]));

	mux_2level_tapbuf_size3 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[90]}),
		.sram(mux_2level_tapbuf_size3_48_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_48_sram_inv[0:1]),
		.out(chany_top_out[60]));

	mux_2level_tapbuf_size3 mux_top_track_122 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[89]}),
		.sram(mux_2level_tapbuf_size3_49_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_49_sram_inv[0:1]),
		.out(chany_top_out[61]));

	mux_2level_tapbuf_size3 mux_top_track_124 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[88]}),
		.sram(mux_2level_tapbuf_size3_50_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_50_sram_inv[0:1]),
		.out(chany_top_out[62]));

	mux_2level_tapbuf_size3 mux_top_track_126 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[87]}),
		.sram(mux_2level_tapbuf_size3_51_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_51_sram_inv[0:1]),
		.out(chany_top_out[63]));

	mux_2level_tapbuf_size3 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[86]}),
		.sram(mux_2level_tapbuf_size3_52_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_52_sram_inv[0:1]),
		.out(chany_top_out[64]));

	mux_2level_tapbuf_size3 mux_top_track_130 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[85]}),
		.sram(mux_2level_tapbuf_size3_53_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_53_sram_inv[0:1]),
		.out(chany_top_out[65]));

	mux_2level_tapbuf_size3 mux_top_track_132 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[84]}),
		.sram(mux_2level_tapbuf_size3_54_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_54_sram_inv[0:1]),
		.out(chany_top_out[66]));

	mux_2level_tapbuf_size3 mux_top_track_134 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[83]}),
		.sram(mux_2level_tapbuf_size3_55_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_55_sram_inv[0:1]),
		.out(chany_top_out[67]));

	mux_2level_tapbuf_size3 mux_top_track_140 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[80]}),
		.sram(mux_2level_tapbuf_size3_56_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_56_sram_inv[0:1]),
		.out(chany_top_out[70]));

	mux_2level_tapbuf_size3 mux_top_track_142 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[79]}),
		.sram(mux_2level_tapbuf_size3_57_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_57_sram_inv[0:1]),
		.out(chany_top_out[71]));

	mux_2level_tapbuf_size3 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[78]}),
		.sram(mux_2level_tapbuf_size3_58_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_58_sram_inv[0:1]),
		.out(chany_top_out[72]));

	mux_2level_tapbuf_size3 mux_top_track_146 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[77]}),
		.sram(mux_2level_tapbuf_size3_59_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_59_sram_inv[0:1]),
		.out(chany_top_out[73]));

	mux_2level_tapbuf_size3 mux_top_track_148 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[76]}),
		.sram(mux_2level_tapbuf_size3_60_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_60_sram_inv[0:1]),
		.out(chany_top_out[74]));

	mux_2level_tapbuf_size3 mux_top_track_150 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[75]}),
		.sram(mux_2level_tapbuf_size3_61_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_61_sram_inv[0:1]),
		.out(chany_top_out[75]));

	mux_2level_tapbuf_size3 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[74]}),
		.sram(mux_2level_tapbuf_size3_62_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_62_sram_inv[0:1]),
		.out(chany_top_out[76]));

	mux_2level_tapbuf_size3 mux_top_track_154 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[73]}),
		.sram(mux_2level_tapbuf_size3_63_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_63_sram_inv[0:1]),
		.out(chany_top_out[77]));

	mux_2level_tapbuf_size3 mux_top_track_160 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[70]}),
		.sram(mux_2level_tapbuf_size3_64_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_64_sram_inv[0:1]),
		.out(chany_top_out[80]));

	mux_2level_tapbuf_size3 mux_top_track_162 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[69]}),
		.sram(mux_2level_tapbuf_size3_65_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_65_sram_inv[0:1]),
		.out(chany_top_out[81]));

	mux_2level_tapbuf_size3 mux_top_track_164 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[68]}),
		.sram(mux_2level_tapbuf_size3_66_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_66_sram_inv[0:1]),
		.out(chany_top_out[82]));

	mux_2level_tapbuf_size3 mux_top_track_166 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[67]}),
		.sram(mux_2level_tapbuf_size3_67_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_67_sram_inv[0:1]),
		.out(chany_top_out[83]));

	mux_2level_tapbuf_size3 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[66]}),
		.sram(mux_2level_tapbuf_size3_68_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_68_sram_inv[0:1]),
		.out(chany_top_out[84]));

	mux_2level_tapbuf_size3 mux_top_track_170 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[65]}),
		.sram(mux_2level_tapbuf_size3_69_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_69_sram_inv[0:1]),
		.out(chany_top_out[85]));

	mux_2level_tapbuf_size3 mux_top_track_172 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[64]}),
		.sram(mux_2level_tapbuf_size3_70_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_70_sram_inv[0:1]),
		.out(chany_top_out[86]));

	mux_2level_tapbuf_size3 mux_top_track_174 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[63]}),
		.sram(mux_2level_tapbuf_size3_71_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_71_sram_inv[0:1]),
		.out(chany_top_out[87]));

	mux_2level_tapbuf_size3 mux_top_track_180 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[60]}),
		.sram(mux_2level_tapbuf_size3_72_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_72_sram_inv[0:1]),
		.out(chany_top_out[90]));

	mux_2level_tapbuf_size3 mux_top_track_182 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[59]}),
		.sram(mux_2level_tapbuf_size3_73_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_73_sram_inv[0:1]),
		.out(chany_top_out[91]));

	mux_2level_tapbuf_size3 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[58]}),
		.sram(mux_2level_tapbuf_size3_74_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_74_sram_inv[0:1]),
		.out(chany_top_out[92]));

	mux_2level_tapbuf_size3 mux_top_track_186 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[57]}),
		.sram(mux_2level_tapbuf_size3_75_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_75_sram_inv[0:1]),
		.out(chany_top_out[93]));

	mux_2level_tapbuf_size3 mux_top_track_188 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[56]}),
		.sram(mux_2level_tapbuf_size3_76_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_76_sram_inv[0:1]),
		.out(chany_top_out[94]));

	mux_2level_tapbuf_size3 mux_top_track_190 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[55]}),
		.sram(mux_2level_tapbuf_size3_77_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_77_sram_inv[0:1]),
		.out(chany_top_out[95]));

	mux_2level_tapbuf_size3 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[54]}),
		.sram(mux_2level_tapbuf_size3_78_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_78_sram_inv[0:1]),
		.out(chany_top_out[96]));

	mux_2level_tapbuf_size3 mux_top_track_194 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[53]}),
		.sram(mux_2level_tapbuf_size3_79_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_79_sram_inv[0:1]),
		.out(chany_top_out[97]));

	mux_2level_tapbuf_size3 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[50]}),
		.sram(mux_2level_tapbuf_size3_80_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_80_sram_inv[0:1]),
		.out(chany_top_out[100]));

	mux_2level_tapbuf_size3 mux_top_track_202 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[49]}),
		.sram(mux_2level_tapbuf_size3_81_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_81_sram_inv[0:1]),
		.out(chany_top_out[101]));

	mux_2level_tapbuf_size3 mux_top_track_204 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[48]}),
		.sram(mux_2level_tapbuf_size3_82_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_82_sram_inv[0:1]),
		.out(chany_top_out[102]));

	mux_2level_tapbuf_size3 mux_top_track_206 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[47]}),
		.sram(mux_2level_tapbuf_size3_83_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_83_sram_inv[0:1]),
		.out(chany_top_out[103]));

	mux_2level_tapbuf_size3 mux_top_track_208 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[46]}),
		.sram(mux_2level_tapbuf_size3_84_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_84_sram_inv[0:1]),
		.out(chany_top_out[104]));

	mux_2level_tapbuf_size3 mux_top_track_210 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[45]}),
		.sram(mux_2level_tapbuf_size3_85_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_85_sram_inv[0:1]),
		.out(chany_top_out[105]));

	mux_2level_tapbuf_size3 mux_top_track_212 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[44]}),
		.sram(mux_2level_tapbuf_size3_86_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_86_sram_inv[0:1]),
		.out(chany_top_out[106]));

	mux_2level_tapbuf_size3 mux_top_track_214 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[43]}),
		.sram(mux_2level_tapbuf_size3_87_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_87_sram_inv[0:1]),
		.out(chany_top_out[107]));

	mux_2level_tapbuf_size3 mux_top_track_220 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[40]}),
		.sram(mux_2level_tapbuf_size3_88_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_88_sram_inv[0:1]),
		.out(chany_top_out[110]));

	mux_2level_tapbuf_size3 mux_top_track_222 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[39]}),
		.sram(mux_2level_tapbuf_size3_89_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_89_sram_inv[0:1]),
		.out(chany_top_out[111]));

	mux_2level_tapbuf_size3 mux_top_track_224 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[38]}),
		.sram(mux_2level_tapbuf_size3_90_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_90_sram_inv[0:1]),
		.out(chany_top_out[112]));

	mux_2level_tapbuf_size3 mux_top_track_226 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[37]}),
		.sram(mux_2level_tapbuf_size3_91_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_91_sram_inv[0:1]),
		.out(chany_top_out[113]));

	mux_2level_tapbuf_size3 mux_top_track_228 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[36]}),
		.sram(mux_2level_tapbuf_size3_92_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_92_sram_inv[0:1]),
		.out(chany_top_out[114]));

	mux_2level_tapbuf_size3 mux_top_track_230 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[35]}),
		.sram(mux_2level_tapbuf_size3_93_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_93_sram_inv[0:1]),
		.out(chany_top_out[115]));

	mux_2level_tapbuf_size3 mux_top_track_232 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[34]}),
		.sram(mux_2level_tapbuf_size3_94_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_94_sram_inv[0:1]),
		.out(chany_top_out[116]));

	mux_2level_tapbuf_size3 mux_top_track_234 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[33]}),
		.sram(mux_2level_tapbuf_size3_95_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_95_sram_inv[0:1]),
		.out(chany_top_out[117]));

	mux_2level_tapbuf_size3 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[30]}),
		.sram(mux_2level_tapbuf_size3_96_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_96_sram_inv[0:1]),
		.out(chany_top_out[120]));

	mux_2level_tapbuf_size3 mux_top_track_242 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[29]}),
		.sram(mux_2level_tapbuf_size3_97_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_97_sram_inv[0:1]),
		.out(chany_top_out[121]));

	mux_2level_tapbuf_size3 mux_top_track_244 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[28]}),
		.sram(mux_2level_tapbuf_size3_98_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_98_sram_inv[0:1]),
		.out(chany_top_out[122]));

	mux_2level_tapbuf_size3 mux_top_track_246 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[27]}),
		.sram(mux_2level_tapbuf_size3_99_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_99_sram_inv[0:1]),
		.out(chany_top_out[123]));

	mux_2level_tapbuf_size3 mux_top_track_248 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[26]}),
		.sram(mux_2level_tapbuf_size3_100_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_100_sram_inv[0:1]),
		.out(chany_top_out[124]));

	mux_2level_tapbuf_size3 mux_top_track_250 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[25]}),
		.sram(mux_2level_tapbuf_size3_101_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_101_sram_inv[0:1]),
		.out(chany_top_out[125]));

	mux_2level_tapbuf_size3 mux_top_track_252 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[24]}),
		.sram(mux_2level_tapbuf_size3_102_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_102_sram_inv[0:1]),
		.out(chany_top_out[126]));

	mux_2level_tapbuf_size3 mux_top_track_254 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[23]}),
		.sram(mux_2level_tapbuf_size3_103_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_103_sram_inv[0:1]),
		.out(chany_top_out[127]));

	mux_2level_tapbuf_size3 mux_top_track_260 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[20]}),
		.sram(mux_2level_tapbuf_size3_104_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_104_sram_inv[0:1]),
		.out(chany_top_out[130]));

	mux_2level_tapbuf_size3 mux_top_track_262 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[19]}),
		.sram(mux_2level_tapbuf_size3_105_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_105_sram_inv[0:1]),
		.out(chany_top_out[131]));

	mux_2level_tapbuf_size3 mux_top_track_264 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[18]}),
		.sram(mux_2level_tapbuf_size3_106_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_106_sram_inv[0:1]),
		.out(chany_top_out[132]));

	mux_2level_tapbuf_size3 mux_top_track_266 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[17]}),
		.sram(mux_2level_tapbuf_size3_107_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_107_sram_inv[0:1]),
		.out(chany_top_out[133]));

	mux_2level_tapbuf_size3 mux_top_track_268 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[16]}),
		.sram(mux_2level_tapbuf_size3_108_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_108_sram_inv[0:1]),
		.out(chany_top_out[134]));

	mux_2level_tapbuf_size3 mux_top_track_270 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[15]}),
		.sram(mux_2level_tapbuf_size3_109_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_109_sram_inv[0:1]),
		.out(chany_top_out[135]));

	mux_2level_tapbuf_size3 mux_top_track_272 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[14]}),
		.sram(mux_2level_tapbuf_size3_110_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_110_sram_inv[0:1]),
		.out(chany_top_out[136]));

	mux_2level_tapbuf_size3 mux_top_track_274 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[13]}),
		.sram(mux_2level_tapbuf_size3_111_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_111_sram_inv[0:1]),
		.out(chany_top_out[137]));

	mux_2level_tapbuf_size3 mux_top_track_280 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[10]}),
		.sram(mux_2level_tapbuf_size3_112_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_112_sram_inv[0:1]),
		.out(chany_top_out[140]));

	mux_2level_tapbuf_size3 mux_top_track_282 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[9]}),
		.sram(mux_2level_tapbuf_size3_113_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_113_sram_inv[0:1]),
		.out(chany_top_out[141]));

	mux_2level_tapbuf_size3 mux_top_track_284 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[8]}),
		.sram(mux_2level_tapbuf_size3_114_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_114_sram_inv[0:1]),
		.out(chany_top_out[142]));

	mux_2level_tapbuf_size3 mux_top_track_286 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[7]}),
		.sram(mux_2level_tapbuf_size3_115_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_115_sram_inv[0:1]),
		.out(chany_top_out[143]));

	mux_2level_tapbuf_size3 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[6]}),
		.sram(mux_2level_tapbuf_size3_116_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_116_sram_inv[0:1]),
		.out(chany_top_out[144]));

	mux_2level_tapbuf_size3 mux_top_track_290 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[5]}),
		.sram(mux_2level_tapbuf_size3_117_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_117_sram_inv[0:1]),
		.out(chany_top_out[145]));

	mux_2level_tapbuf_size3 mux_top_track_292 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[4]}),
		.sram(mux_2level_tapbuf_size3_118_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_118_sram_inv[0:1]),
		.out(chany_top_out[146]));

	mux_2level_tapbuf_size3 mux_top_track_294 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[3]}),
		.sram(mux_2level_tapbuf_size3_119_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_119_sram_inv[0:1]),
		.out(chany_top_out[147]));

	mux_2level_tapbuf_size3 mux_left_track_1 (
		.in({chany_top_in[0], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_120_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_120_sram_inv[0:1]),
		.out(chanx_left_out[0]));

	mux_2level_tapbuf_size3 mux_left_track_3 (
		.in({chany_top_in[149], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_121_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_121_sram_inv[0:1]),
		.out(chanx_left_out[1]));

	mux_2level_tapbuf_size3 mux_left_track_5 (
		.in({chany_top_in[148], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_122_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_122_sram_inv[0:1]),
		.out(chanx_left_out[2]));

	mux_2level_tapbuf_size3 mux_left_track_7 (
		.in({chany_top_in[147], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_123_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_123_sram_inv[0:1]),
		.out(chanx_left_out[3]));

	mux_2level_tapbuf_size3 mux_left_track_9 (
		.in({chany_top_in[146], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_124_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_124_sram_inv[0:1]),
		.out(chanx_left_out[4]));

	mux_2level_tapbuf_size3 mux_left_track_11 (
		.in({chany_top_in[145], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_125_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_125_sram_inv[0:1]),
		.out(chanx_left_out[5]));

	mux_2level_tapbuf_size3 mux_left_track_13 (
		.in({chany_top_in[144], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_126_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_126_sram_inv[0:1]),
		.out(chanx_left_out[6]));

	mux_2level_tapbuf_size3 mux_left_track_15 (
		.in({chany_top_in[143], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_127_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_127_sram_inv[0:1]),
		.out(chanx_left_out[7]));

	mux_2level_tapbuf_size3 mux_left_track_21 (
		.in({chany_top_in[140], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_128_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_128_sram_inv[0:1]),
		.out(chanx_left_out[10]));

	mux_2level_tapbuf_size3 mux_left_track_23 (
		.in({chany_top_in[139], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_129_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_129_sram_inv[0:1]),
		.out(chanx_left_out[11]));

	mux_2level_tapbuf_size3 mux_left_track_25 (
		.in({chany_top_in[138], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_130_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_130_sram_inv[0:1]),
		.out(chanx_left_out[12]));

	mux_2level_tapbuf_size3 mux_left_track_27 (
		.in({chany_top_in[137], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_131_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_131_sram_inv[0:1]),
		.out(chanx_left_out[13]));

	mux_2level_tapbuf_size3 mux_left_track_29 (
		.in({chany_top_in[136], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_132_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_132_sram_inv[0:1]),
		.out(chanx_left_out[14]));

	mux_2level_tapbuf_size3 mux_left_track_31 (
		.in({chany_top_in[135], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_133_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_133_sram_inv[0:1]),
		.out(chanx_left_out[15]));

	mux_2level_tapbuf_size3 mux_left_track_33 (
		.in({chany_top_in[134], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_134_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_134_sram_inv[0:1]),
		.out(chanx_left_out[16]));

	mux_2level_tapbuf_size3 mux_left_track_35 (
		.in({chany_top_in[133], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_135_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_135_sram_inv[0:1]),
		.out(chanx_left_out[17]));

	mux_2level_tapbuf_size3 mux_left_track_41 (
		.in({chany_top_in[130], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_136_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_136_sram_inv[0:1]),
		.out(chanx_left_out[20]));

	mux_2level_tapbuf_size3 mux_left_track_43 (
		.in({chany_top_in[129], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_137_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_137_sram_inv[0:1]),
		.out(chanx_left_out[21]));

	mux_2level_tapbuf_size3 mux_left_track_45 (
		.in({chany_top_in[128], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_138_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_138_sram_inv[0:1]),
		.out(chanx_left_out[22]));

	mux_2level_tapbuf_size3 mux_left_track_47 (
		.in({chany_top_in[127], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_139_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_139_sram_inv[0:1]),
		.out(chanx_left_out[23]));

	mux_2level_tapbuf_size3 mux_left_track_49 (
		.in({chany_top_in[126], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_140_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_140_sram_inv[0:1]),
		.out(chanx_left_out[24]));

	mux_2level_tapbuf_size3 mux_left_track_51 (
		.in({chany_top_in[125], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_141_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_141_sram_inv[0:1]),
		.out(chanx_left_out[25]));

	mux_2level_tapbuf_size3 mux_left_track_53 (
		.in({chany_top_in[124], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_142_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_142_sram_inv[0:1]),
		.out(chanx_left_out[26]));

	mux_2level_tapbuf_size3 mux_left_track_55 (
		.in({chany_top_in[123], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_143_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_143_sram_inv[0:1]),
		.out(chanx_left_out[27]));

	mux_2level_tapbuf_size3 mux_left_track_61 (
		.in({chany_top_in[120], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_144_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_144_sram_inv[0:1]),
		.out(chanx_left_out[30]));

	mux_2level_tapbuf_size3 mux_left_track_63 (
		.in({chany_top_in[119], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_145_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_145_sram_inv[0:1]),
		.out(chanx_left_out[31]));

	mux_2level_tapbuf_size3 mux_left_track_65 (
		.in({chany_top_in[118], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_146_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_146_sram_inv[0:1]),
		.out(chanx_left_out[32]));

	mux_2level_tapbuf_size3 mux_left_track_67 (
		.in({chany_top_in[117], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_147_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_147_sram_inv[0:1]),
		.out(chanx_left_out[33]));

	mux_2level_tapbuf_size3 mux_left_track_69 (
		.in({chany_top_in[116], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_148_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_148_sram_inv[0:1]),
		.out(chanx_left_out[34]));

	mux_2level_tapbuf_size3 mux_left_track_71 (
		.in({chany_top_in[115], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_149_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_149_sram_inv[0:1]),
		.out(chanx_left_out[35]));

	mux_2level_tapbuf_size3 mux_left_track_73 (
		.in({chany_top_in[114], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_150_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_150_sram_inv[0:1]),
		.out(chanx_left_out[36]));

	mux_2level_tapbuf_size3 mux_left_track_75 (
		.in({chany_top_in[113], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_151_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_151_sram_inv[0:1]),
		.out(chanx_left_out[37]));

	mux_2level_tapbuf_size3 mux_left_track_81 (
		.in({chany_top_in[110], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_152_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_152_sram_inv[0:1]),
		.out(chanx_left_out[40]));

	mux_2level_tapbuf_size3 mux_left_track_83 (
		.in({chany_top_in[109], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_153_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_153_sram_inv[0:1]),
		.out(chanx_left_out[41]));

	mux_2level_tapbuf_size3 mux_left_track_85 (
		.in({chany_top_in[108], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_154_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_154_sram_inv[0:1]),
		.out(chanx_left_out[42]));

	mux_2level_tapbuf_size3 mux_left_track_87 (
		.in({chany_top_in[107], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_155_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_155_sram_inv[0:1]),
		.out(chanx_left_out[43]));

	mux_2level_tapbuf_size3 mux_left_track_89 (
		.in({chany_top_in[106], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_156_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_156_sram_inv[0:1]),
		.out(chanx_left_out[44]));

	mux_2level_tapbuf_size3 mux_left_track_91 (
		.in({chany_top_in[105], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_157_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_157_sram_inv[0:1]),
		.out(chanx_left_out[45]));

	mux_2level_tapbuf_size3 mux_left_track_93 (
		.in({chany_top_in[104], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_158_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_158_sram_inv[0:1]),
		.out(chanx_left_out[46]));

	mux_2level_tapbuf_size3 mux_left_track_95 (
		.in({chany_top_in[103], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_159_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_159_sram_inv[0:1]),
		.out(chanx_left_out[47]));

	mux_2level_tapbuf_size3 mux_left_track_101 (
		.in({chany_top_in[100], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_160_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_160_sram_inv[0:1]),
		.out(chanx_left_out[50]));

	mux_2level_tapbuf_size3 mux_left_track_103 (
		.in({chany_top_in[99], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_161_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_161_sram_inv[0:1]),
		.out(chanx_left_out[51]));

	mux_2level_tapbuf_size3 mux_left_track_105 (
		.in({chany_top_in[98], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_162_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_162_sram_inv[0:1]),
		.out(chanx_left_out[52]));

	mux_2level_tapbuf_size3 mux_left_track_107 (
		.in({chany_top_in[97], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_163_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_163_sram_inv[0:1]),
		.out(chanx_left_out[53]));

	mux_2level_tapbuf_size3 mux_left_track_109 (
		.in({chany_top_in[96], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_164_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_164_sram_inv[0:1]),
		.out(chanx_left_out[54]));

	mux_2level_tapbuf_size3 mux_left_track_111 (
		.in({chany_top_in[95], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_165_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_165_sram_inv[0:1]),
		.out(chanx_left_out[55]));

	mux_2level_tapbuf_size3 mux_left_track_113 (
		.in({chany_top_in[94], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_166_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_166_sram_inv[0:1]),
		.out(chanx_left_out[56]));

	mux_2level_tapbuf_size3 mux_left_track_115 (
		.in({chany_top_in[93], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_167_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_167_sram_inv[0:1]),
		.out(chanx_left_out[57]));

	mux_2level_tapbuf_size3 mux_left_track_121 (
		.in({chany_top_in[90], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_168_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_168_sram_inv[0:1]),
		.out(chanx_left_out[60]));

	mux_2level_tapbuf_size3 mux_left_track_123 (
		.in({chany_top_in[89], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_169_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_169_sram_inv[0:1]),
		.out(chanx_left_out[61]));

	mux_2level_tapbuf_size3 mux_left_track_125 (
		.in({chany_top_in[88], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_170_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_170_sram_inv[0:1]),
		.out(chanx_left_out[62]));

	mux_2level_tapbuf_size3 mux_left_track_127 (
		.in({chany_top_in[87], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_171_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_171_sram_inv[0:1]),
		.out(chanx_left_out[63]));

	mux_2level_tapbuf_size3 mux_left_track_129 (
		.in({chany_top_in[86], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_172_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_172_sram_inv[0:1]),
		.out(chanx_left_out[64]));

	mux_2level_tapbuf_size3 mux_left_track_131 (
		.in({chany_top_in[85], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_173_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_173_sram_inv[0:1]),
		.out(chanx_left_out[65]));

	mux_2level_tapbuf_size3 mux_left_track_133 (
		.in({chany_top_in[84], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_174_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_174_sram_inv[0:1]),
		.out(chanx_left_out[66]));

	mux_2level_tapbuf_size3 mux_left_track_135 (
		.in({chany_top_in[83], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_175_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_175_sram_inv[0:1]),
		.out(chanx_left_out[67]));

	mux_2level_tapbuf_size3 mux_left_track_141 (
		.in({chany_top_in[80], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_176_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_176_sram_inv[0:1]),
		.out(chanx_left_out[70]));

	mux_2level_tapbuf_size3 mux_left_track_143 (
		.in({chany_top_in[79], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_177_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_177_sram_inv[0:1]),
		.out(chanx_left_out[71]));

	mux_2level_tapbuf_size3 mux_left_track_145 (
		.in({chany_top_in[78], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_178_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_178_sram_inv[0:1]),
		.out(chanx_left_out[72]));

	mux_2level_tapbuf_size3 mux_left_track_147 (
		.in({chany_top_in[77], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_179_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_179_sram_inv[0:1]),
		.out(chanx_left_out[73]));

	mux_2level_tapbuf_size3 mux_left_track_149 (
		.in({chany_top_in[76], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_180_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_180_sram_inv[0:1]),
		.out(chanx_left_out[74]));

	mux_2level_tapbuf_size3 mux_left_track_151 (
		.in({chany_top_in[75], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_181_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_181_sram_inv[0:1]),
		.out(chanx_left_out[75]));

	mux_2level_tapbuf_size3 mux_left_track_153 (
		.in({chany_top_in[74], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_182_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_182_sram_inv[0:1]),
		.out(chanx_left_out[76]));

	mux_2level_tapbuf_size3 mux_left_track_155 (
		.in({chany_top_in[73], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_183_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_183_sram_inv[0:1]),
		.out(chanx_left_out[77]));

	mux_2level_tapbuf_size3 mux_left_track_161 (
		.in({chany_top_in[70], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_184_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_184_sram_inv[0:1]),
		.out(chanx_left_out[80]));

	mux_2level_tapbuf_size3 mux_left_track_163 (
		.in({chany_top_in[69], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_185_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_185_sram_inv[0:1]),
		.out(chanx_left_out[81]));

	mux_2level_tapbuf_size3 mux_left_track_165 (
		.in({chany_top_in[68], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_186_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_186_sram_inv[0:1]),
		.out(chanx_left_out[82]));

	mux_2level_tapbuf_size3 mux_left_track_167 (
		.in({chany_top_in[67], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_187_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_187_sram_inv[0:1]),
		.out(chanx_left_out[83]));

	mux_2level_tapbuf_size3 mux_left_track_169 (
		.in({chany_top_in[66], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_188_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_188_sram_inv[0:1]),
		.out(chanx_left_out[84]));

	mux_2level_tapbuf_size3 mux_left_track_171 (
		.in({chany_top_in[65], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_189_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_189_sram_inv[0:1]),
		.out(chanx_left_out[85]));

	mux_2level_tapbuf_size3 mux_left_track_173 (
		.in({chany_top_in[64], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_190_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_190_sram_inv[0:1]),
		.out(chanx_left_out[86]));

	mux_2level_tapbuf_size3 mux_left_track_175 (
		.in({chany_top_in[63], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_191_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_191_sram_inv[0:1]),
		.out(chanx_left_out[87]));

	mux_2level_tapbuf_size3 mux_left_track_181 (
		.in({chany_top_in[60], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_192_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_192_sram_inv[0:1]),
		.out(chanx_left_out[90]));

	mux_2level_tapbuf_size3 mux_left_track_183 (
		.in({chany_top_in[59], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_193_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_193_sram_inv[0:1]),
		.out(chanx_left_out[91]));

	mux_2level_tapbuf_size3 mux_left_track_185 (
		.in({chany_top_in[58], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_194_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_194_sram_inv[0:1]),
		.out(chanx_left_out[92]));

	mux_2level_tapbuf_size3 mux_left_track_187 (
		.in({chany_top_in[57], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_195_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_195_sram_inv[0:1]),
		.out(chanx_left_out[93]));

	mux_2level_tapbuf_size3 mux_left_track_189 (
		.in({chany_top_in[56], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_196_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_196_sram_inv[0:1]),
		.out(chanx_left_out[94]));

	mux_2level_tapbuf_size3 mux_left_track_191 (
		.in({chany_top_in[55], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_197_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_197_sram_inv[0:1]),
		.out(chanx_left_out[95]));

	mux_2level_tapbuf_size3 mux_left_track_193 (
		.in({chany_top_in[54], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_198_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_198_sram_inv[0:1]),
		.out(chanx_left_out[96]));

	mux_2level_tapbuf_size3 mux_left_track_195 (
		.in({chany_top_in[53], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_199_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_199_sram_inv[0:1]),
		.out(chanx_left_out[97]));

	mux_2level_tapbuf_size3 mux_left_track_201 (
		.in({chany_top_in[50], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_200_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_200_sram_inv[0:1]),
		.out(chanx_left_out[100]));

	mux_2level_tapbuf_size3 mux_left_track_203 (
		.in({chany_top_in[49], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_201_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_201_sram_inv[0:1]),
		.out(chanx_left_out[101]));

	mux_2level_tapbuf_size3 mux_left_track_205 (
		.in({chany_top_in[48], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_202_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_202_sram_inv[0:1]),
		.out(chanx_left_out[102]));

	mux_2level_tapbuf_size3 mux_left_track_207 (
		.in({chany_top_in[47], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_203_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_203_sram_inv[0:1]),
		.out(chanx_left_out[103]));

	mux_2level_tapbuf_size3 mux_left_track_209 (
		.in({chany_top_in[46], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_204_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_204_sram_inv[0:1]),
		.out(chanx_left_out[104]));

	mux_2level_tapbuf_size3 mux_left_track_211 (
		.in({chany_top_in[45], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_205_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_205_sram_inv[0:1]),
		.out(chanx_left_out[105]));

	mux_2level_tapbuf_size3 mux_left_track_213 (
		.in({chany_top_in[44], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_206_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_206_sram_inv[0:1]),
		.out(chanx_left_out[106]));

	mux_2level_tapbuf_size3 mux_left_track_215 (
		.in({chany_top_in[43], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_207_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_207_sram_inv[0:1]),
		.out(chanx_left_out[107]));

	mux_2level_tapbuf_size3 mux_left_track_221 (
		.in({chany_top_in[40], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_208_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_208_sram_inv[0:1]),
		.out(chanx_left_out[110]));

	mux_2level_tapbuf_size3 mux_left_track_223 (
		.in({chany_top_in[39], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_209_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_209_sram_inv[0:1]),
		.out(chanx_left_out[111]));

	mux_2level_tapbuf_size3 mux_left_track_225 (
		.in({chany_top_in[38], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_210_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_210_sram_inv[0:1]),
		.out(chanx_left_out[112]));

	mux_2level_tapbuf_size3 mux_left_track_227 (
		.in({chany_top_in[37], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_211_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_211_sram_inv[0:1]),
		.out(chanx_left_out[113]));

	mux_2level_tapbuf_size3 mux_left_track_229 (
		.in({chany_top_in[36], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_212_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_212_sram_inv[0:1]),
		.out(chanx_left_out[114]));

	mux_2level_tapbuf_size3 mux_left_track_231 (
		.in({chany_top_in[35], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_213_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_213_sram_inv[0:1]),
		.out(chanx_left_out[115]));

	mux_2level_tapbuf_size3 mux_left_track_233 (
		.in({chany_top_in[34], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_214_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_214_sram_inv[0:1]),
		.out(chanx_left_out[116]));

	mux_2level_tapbuf_size3 mux_left_track_235 (
		.in({chany_top_in[33], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_215_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_215_sram_inv[0:1]),
		.out(chanx_left_out[117]));

	mux_2level_tapbuf_size3 mux_left_track_241 (
		.in({chany_top_in[30], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_216_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_216_sram_inv[0:1]),
		.out(chanx_left_out[120]));

	mux_2level_tapbuf_size3 mux_left_track_243 (
		.in({chany_top_in[29], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_217_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_217_sram_inv[0:1]),
		.out(chanx_left_out[121]));

	mux_2level_tapbuf_size3 mux_left_track_245 (
		.in({chany_top_in[28], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_218_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_218_sram_inv[0:1]),
		.out(chanx_left_out[122]));

	mux_2level_tapbuf_size3 mux_left_track_247 (
		.in({chany_top_in[27], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_219_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_219_sram_inv[0:1]),
		.out(chanx_left_out[123]));

	mux_2level_tapbuf_size3 mux_left_track_249 (
		.in({chany_top_in[26], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_220_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_220_sram_inv[0:1]),
		.out(chanx_left_out[124]));

	mux_2level_tapbuf_size3 mux_left_track_251 (
		.in({chany_top_in[25], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_221_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_221_sram_inv[0:1]),
		.out(chanx_left_out[125]));

	mux_2level_tapbuf_size3 mux_left_track_253 (
		.in({chany_top_in[24], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_222_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_222_sram_inv[0:1]),
		.out(chanx_left_out[126]));

	mux_2level_tapbuf_size3 mux_left_track_255 (
		.in({chany_top_in[23], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_223_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_223_sram_inv[0:1]),
		.out(chanx_left_out[127]));

	mux_2level_tapbuf_size3 mux_left_track_261 (
		.in({chany_top_in[20], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_224_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_224_sram_inv[0:1]),
		.out(chanx_left_out[130]));

	mux_2level_tapbuf_size3 mux_left_track_263 (
		.in({chany_top_in[19], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_225_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_225_sram_inv[0:1]),
		.out(chanx_left_out[131]));

	mux_2level_tapbuf_size3 mux_left_track_265 (
		.in({chany_top_in[18], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_226_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_226_sram_inv[0:1]),
		.out(chanx_left_out[132]));

	mux_2level_tapbuf_size3 mux_left_track_267 (
		.in({chany_top_in[17], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_227_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_227_sram_inv[0:1]),
		.out(chanx_left_out[133]));

	mux_2level_tapbuf_size3 mux_left_track_269 (
		.in({chany_top_in[16], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_228_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_228_sram_inv[0:1]),
		.out(chanx_left_out[134]));

	mux_2level_tapbuf_size3 mux_left_track_271 (
		.in({chany_top_in[15], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_229_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_229_sram_inv[0:1]),
		.out(chanx_left_out[135]));

	mux_2level_tapbuf_size3 mux_left_track_273 (
		.in({chany_top_in[14], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_230_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_230_sram_inv[0:1]),
		.out(chanx_left_out[136]));

	mux_2level_tapbuf_size3 mux_left_track_275 (
		.in({chany_top_in[13], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_231_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_231_sram_inv[0:1]),
		.out(chanx_left_out[137]));

	mux_2level_tapbuf_size3 mux_left_track_281 (
		.in({chany_top_in[10], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_232_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_232_sram_inv[0:1]),
		.out(chanx_left_out[140]));

	mux_2level_tapbuf_size3 mux_left_track_283 (
		.in({chany_top_in[9], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_233_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_233_sram_inv[0:1]),
		.out(chanx_left_out[141]));

	mux_2level_tapbuf_size3 mux_left_track_285 (
		.in({chany_top_in[8], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_234_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_234_sram_inv[0:1]),
		.out(chanx_left_out[142]));

	mux_2level_tapbuf_size3 mux_left_track_287 (
		.in({chany_top_in[7], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_235_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_235_sram_inv[0:1]),
		.out(chanx_left_out[143]));

	mux_2level_tapbuf_size3 mux_left_track_289 (
		.in({chany_top_in[6], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_236_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_236_sram_inv[0:1]),
		.out(chanx_left_out[144]));

	mux_2level_tapbuf_size3 mux_left_track_291 (
		.in({chany_top_in[5], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_237_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_237_sram_inv[0:1]),
		.out(chanx_left_out[145]));

	mux_2level_tapbuf_size3 mux_left_track_293 (
		.in({chany_top_in[4], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_238_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_238_sram_inv[0:1]),
		.out(chanx_left_out[146]));

	mux_2level_tapbuf_size3 mux_left_track_295 (
		.in({chany_top_in[3], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_239_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_239_sram_inv[0:1]),
		.out(chanx_left_out[147]));

	mux_2level_tapbuf_size3_mem mem_top_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_0_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_1_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_2_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_6 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_3_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_4_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_5_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_6_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_14 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_7_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_8_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_22 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_9_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_10_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_11_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_12_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_30 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_13_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_14_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_34 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_15_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_16_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_17_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_18_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_46 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_19_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_20_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_21_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_52 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_22_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_54 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_23_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_24_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_62 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_25_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_26_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_27_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_28_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_70 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_29_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_30_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_31_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_32_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_33_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_33_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_34_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_34_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_86 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_35_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_35_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_36_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_36_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_37_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_37_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_38_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_38_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_94 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_39_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_39_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_40_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_40_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_102 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_41_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_41_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_42_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_42_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_106 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_43_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_43_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_44_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_44_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_110 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_45_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_45_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_46_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_46_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_47_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_47_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_48_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_48_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_49_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_49_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_124 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_50_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_50_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_126 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_51_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_51_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_52_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_52_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_53_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_53_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_54_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_54_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_134 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_55_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_55_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_56_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_56_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_142 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_57_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_57_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_58_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_58_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_59_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_59_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_60_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_60_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_150 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_61_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_61_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_62_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_62_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_63_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_63_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_64_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_64_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_65_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_65_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_66_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_66_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_166 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_67_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_67_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_68_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_68_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_69_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_69_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_70_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_70_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_174 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_71_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_71_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_72_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_72_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_182 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_73_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_73_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_74_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_74_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_75_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_75_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_76_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_76_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_190 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_77_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_77_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_78_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_78_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_78_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_79_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_79_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_79_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_80_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_80_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_80_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_80_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_81_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_81_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_81_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_81_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_82_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_82_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_82_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_206 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_82_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_83_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_83_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_83_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_83_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_84_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_84_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_84_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_210 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_84_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_85_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_85_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_85_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_212 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_85_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_86_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_86_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_86_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_214 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_86_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_87_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_87_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_87_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_220 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_88_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_88_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_88_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_222 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_88_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_89_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_89_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_89_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_89_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_90_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_90_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_90_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_226 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_90_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_91_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_91_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_91_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_228 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_91_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_92_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_92_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_92_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_230 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_92_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_93_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_93_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_93_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_93_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_94_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_94_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_94_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_234 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_94_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_95_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_95_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_95_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_96_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_96_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_96_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_242 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_96_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_97_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_97_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_97_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_244 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_97_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_98_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_98_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_98_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_246 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_98_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_99_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_99_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_99_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_99_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_100_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_100_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_100_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_250 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_100_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_101_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_101_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_101_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_252 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_101_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_102_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_102_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_102_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_254 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_102_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_103_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_103_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_103_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_260 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_104_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_104_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_104_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_262 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_104_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_105_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_105_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_105_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_105_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_106_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_106_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_106_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_266 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_106_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_107_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_107_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_107_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_268 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_107_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_108_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_108_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_108_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_270 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_108_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_109_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_109_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_109_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_109_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_110_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_110_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_110_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_274 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_110_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_111_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_111_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_111_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_112_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_112_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_112_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_282 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_112_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_113_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_113_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_113_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_284 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_113_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_114_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_114_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_114_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_286 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_114_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_115_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_115_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_115_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_115_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_116_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_116_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_116_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_290 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_116_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_117_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_117_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_117_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_292 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_117_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_118_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_118_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_118_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_294 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_118_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_119_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_119_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_119_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_120_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_120_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_120_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_3 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_120_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_121_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_121_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_121_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_5 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_121_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_122_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_122_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_122_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_7 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_122_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_123_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_123_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_123_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_123_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_124_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_124_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_124_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_11 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_124_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_125_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_125_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_125_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_13 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_125_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_126_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_126_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_126_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_15 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_126_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_127_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_127_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_127_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_21 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_128_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_128_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_128_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_23 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_128_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_129_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_129_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_129_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_129_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_130_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_130_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_130_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_27 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_130_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_131_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_131_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_131_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_29 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_131_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_132_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_132_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_132_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_31 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_132_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_133_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_133_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_133_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_133_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_134_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_134_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_134_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_35 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_134_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_135_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_135_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_135_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_136_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_136_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_136_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_43 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_136_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_137_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_137_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_137_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_45 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_137_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_138_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_138_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_138_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_47 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_138_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_139_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_139_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_139_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_139_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_140_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_140_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_140_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_51 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_140_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_141_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_141_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_141_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_53 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_141_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_142_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_142_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_142_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_55 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_142_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_143_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_143_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_143_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_61 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_144_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_144_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_144_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_63 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_144_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_145_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_145_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_145_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_145_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_146_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_146_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_146_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_67 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_146_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_147_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_147_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_147_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_69 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_147_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_148_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_148_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_148_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_71 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_148_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_149_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_149_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_149_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_149_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_150_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_150_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_150_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_75 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_150_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_151_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_151_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_151_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_152_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_152_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_152_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_83 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_152_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_153_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_153_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_153_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_85 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_153_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_154_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_154_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_154_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_87 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_154_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_155_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_155_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_155_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_155_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_156_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_156_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_156_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_91 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_156_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_157_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_157_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_157_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_93 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_157_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_158_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_158_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_158_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_95 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_158_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_159_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_159_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_159_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_101 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_160_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_160_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_160_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_103 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_160_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_161_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_161_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_161_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_105 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_161_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_162_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_162_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_162_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_107 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_162_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_163_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_163_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_163_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_109 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_163_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_164_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_164_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_164_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_111 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_164_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_165_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_165_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_165_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_113 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_165_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_166_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_166_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_166_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_115 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_166_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_167_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_167_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_167_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_121 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_168_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_168_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_168_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_123 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_168_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_169_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_169_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_169_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_125 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_169_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_170_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_170_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_170_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_127 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_170_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_171_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_171_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_171_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_129 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_171_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_172_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_172_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_172_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_131 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_172_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_173_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_173_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_173_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_133 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_173_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_174_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_174_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_174_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_135 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_174_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_175_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_175_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_175_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_141 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_176_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_176_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_176_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_143 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_176_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_177_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_177_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_177_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_145 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_177_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_178_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_178_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_178_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_147 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_178_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_179_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_179_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_179_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_149 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_179_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_180_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_180_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_180_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_151 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_180_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_181_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_181_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_181_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_153 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_181_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_182_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_182_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_182_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_155 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_182_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_183_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_183_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_183_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_161 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_184_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_184_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_184_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_163 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_184_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_185_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_185_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_185_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_165 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_185_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_186_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_186_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_186_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_167 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_186_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_187_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_187_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_187_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_169 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_187_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_188_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_188_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_188_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_171 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_188_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_189_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_189_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_189_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_173 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_189_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_190_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_190_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_190_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_175 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_190_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_191_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_191_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_191_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_181 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_192_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_192_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_192_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_183 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_192_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_193_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_193_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_193_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_185 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_193_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_194_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_194_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_194_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_187 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_194_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_195_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_195_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_195_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_189 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_195_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_196_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_196_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_196_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_191 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_196_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_197_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_197_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_197_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_193 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_197_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_198_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_198_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_198_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_195 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_198_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_199_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_199_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_199_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_201 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_200_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_200_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_200_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_203 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_200_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_201_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_201_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_201_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_205 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_201_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_202_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_202_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_202_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_207 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_202_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_203_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_203_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_203_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_209 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_203_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_204_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_204_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_204_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_211 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_204_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_205_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_205_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_205_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_213 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_205_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_206_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_206_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_206_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_215 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_206_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_207_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_207_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_207_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_221 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_208_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_208_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_208_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_223 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_208_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_209_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_209_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_209_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_225 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_209_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_210_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_210_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_210_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_227 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_210_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_211_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_211_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_211_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_229 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_211_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_212_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_212_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_212_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_231 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_212_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_213_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_213_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_213_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_233 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_213_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_214_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_214_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_214_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_235 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_214_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_215_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_215_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_215_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_241 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_216_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_216_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_216_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_243 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_216_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_217_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_217_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_217_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_245 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_217_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_218_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_218_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_218_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_247 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_218_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_219_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_219_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_219_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_249 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_219_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_220_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_220_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_220_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_251 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_220_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_221_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_221_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_221_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_253 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_221_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_222_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_222_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_222_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_255 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_222_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_223_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_223_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_223_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_261 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_224_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_224_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_224_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_263 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_224_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_225_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_225_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_225_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_265 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_225_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_226_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_226_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_226_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_267 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_226_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_227_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_227_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_227_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_269 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_227_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_228_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_228_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_228_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_271 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_228_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_229_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_229_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_229_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_273 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_229_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_230_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_230_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_230_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_275 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_230_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_231_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_231_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_231_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_281 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_232_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_232_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_232_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_283 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_232_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_233_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_233_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_233_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_285 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_233_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_234_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_234_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_234_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_287 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_234_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_235_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_235_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_235_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_289 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_235_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_236_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_236_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_236_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_291 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_236_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_237_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_237_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_237_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_293 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_237_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_238_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_238_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_238_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_left_track_295 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_238_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_239_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_239_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_239_sram_inv[0:1]));

	mux_2level_tapbuf_size2 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[142]}),
		.sram(mux_2level_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_0_sram_inv[0:1]),
		.out(chany_top_out[8]));

	mux_2level_tapbuf_size2 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[141]}),
		.sram(mux_2level_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_1_sram_inv[0:1]),
		.out(chany_top_out[9]));

	mux_2level_tapbuf_size2 mux_top_track_36 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[132]}),
		.sram(mux_2level_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_2_sram_inv[0:1]),
		.out(chany_top_out[18]));

	mux_2level_tapbuf_size2 mux_top_track_38 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[131]}),
		.sram(mux_2level_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_3_sram_inv[0:1]),
		.out(chany_top_out[19]));

	mux_2level_tapbuf_size2 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[122]}),
		.sram(mux_2level_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_4_sram_inv[0:1]),
		.out(chany_top_out[28]));

	mux_2level_tapbuf_size2 mux_top_track_58 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[121]}),
		.sram(mux_2level_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_5_sram_inv[0:1]),
		.out(chany_top_out[29]));

	mux_2level_tapbuf_size2 mux_top_track_76 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[112]}),
		.sram(mux_2level_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_6_sram_inv[0:1]),
		.out(chany_top_out[38]));

	mux_2level_tapbuf_size2 mux_top_track_78 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[111]}),
		.sram(mux_2level_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_7_sram_inv[0:1]),
		.out(chany_top_out[39]));

	mux_2level_tapbuf_size2 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[102]}),
		.sram(mux_2level_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_8_sram_inv[0:1]),
		.out(chany_top_out[48]));

	mux_2level_tapbuf_size2 mux_top_track_98 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[101]}),
		.sram(mux_2level_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_9_sram_inv[0:1]),
		.out(chany_top_out[49]));

	mux_2level_tapbuf_size2 mux_top_track_116 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[92]}),
		.sram(mux_2level_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_10_sram_inv[0:1]),
		.out(chany_top_out[58]));

	mux_2level_tapbuf_size2 mux_top_track_118 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[91]}),
		.sram(mux_2level_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_11_sram_inv[0:1]),
		.out(chany_top_out[59]));

	mux_2level_tapbuf_size2 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[82]}),
		.sram(mux_2level_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_12_sram_inv[0:1]),
		.out(chany_top_out[68]));

	mux_2level_tapbuf_size2 mux_top_track_138 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[81]}),
		.sram(mux_2level_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_13_sram_inv[0:1]),
		.out(chany_top_out[69]));

	mux_2level_tapbuf_size2 mux_top_track_156 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[72]}),
		.sram(mux_2level_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_14_sram_inv[0:1]),
		.out(chany_top_out[78]));

	mux_2level_tapbuf_size2 mux_top_track_158 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[71]}),
		.sram(mux_2level_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_15_sram_inv[0:1]),
		.out(chany_top_out[79]));

	mux_2level_tapbuf_size2 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[62]}),
		.sram(mux_2level_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_16_sram_inv[0:1]),
		.out(chany_top_out[88]));

	mux_2level_tapbuf_size2 mux_top_track_178 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[61]}),
		.sram(mux_2level_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_17_sram_inv[0:1]),
		.out(chany_top_out[89]));

	mux_2level_tapbuf_size2 mux_top_track_196 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[52]}),
		.sram(mux_2level_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_18_sram_inv[0:1]),
		.out(chany_top_out[98]));

	mux_2level_tapbuf_size2 mux_top_track_198 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[51]}),
		.sram(mux_2level_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_19_sram_inv[0:1]),
		.out(chany_top_out[99]));

	mux_2level_tapbuf_size2 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[42]}),
		.sram(mux_2level_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_20_sram_inv[0:1]),
		.out(chany_top_out[108]));

	mux_2level_tapbuf_size2 mux_top_track_218 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[41]}),
		.sram(mux_2level_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_21_sram_inv[0:1]),
		.out(chany_top_out[109]));

	mux_2level_tapbuf_size2 mux_top_track_236 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[32]}),
		.sram(mux_2level_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_22_sram_inv[0:1]),
		.out(chany_top_out[118]));

	mux_2level_tapbuf_size2 mux_top_track_238 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[31]}),
		.sram(mux_2level_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_23_sram_inv[0:1]),
		.out(chany_top_out[119]));

	mux_2level_tapbuf_size2 mux_top_track_256 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[22]}),
		.sram(mux_2level_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_24_sram_inv[0:1]),
		.out(chany_top_out[128]));

	mux_2level_tapbuf_size2 mux_top_track_258 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[21]}),
		.sram(mux_2level_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_25_sram_inv[0:1]),
		.out(chany_top_out[129]));

	mux_2level_tapbuf_size2 mux_top_track_276 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[12]}),
		.sram(mux_2level_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_26_sram_inv[0:1]),
		.out(chany_top_out[138]));

	mux_2level_tapbuf_size2 mux_top_track_278 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[11]}),
		.sram(mux_2level_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_27_sram_inv[0:1]),
		.out(chany_top_out[139]));

	mux_2level_tapbuf_size2 mux_top_track_296 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[2]}),
		.sram(mux_2level_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_28_sram_inv[0:1]),
		.out(chany_top_out[148]));

	mux_2level_tapbuf_size2 mux_top_track_298 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[1]}),
		.sram(mux_2level_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_29_sram_inv[0:1]),
		.out(chany_top_out[149]));

	mux_2level_tapbuf_size2 mux_left_track_17 (
		.in({chany_top_in[142], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_30_sram_inv[0:1]),
		.out(chanx_left_out[8]));

	mux_2level_tapbuf_size2 mux_left_track_19 (
		.in({chany_top_in[141], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_31_sram_inv[0:1]),
		.out(chanx_left_out[9]));

	mux_2level_tapbuf_size2 mux_left_track_37 (
		.in({chany_top_in[132], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_32_sram_inv[0:1]),
		.out(chanx_left_out[18]));

	mux_2level_tapbuf_size2 mux_left_track_39 (
		.in({chany_top_in[131], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_33_sram_inv[0:1]),
		.out(chanx_left_out[19]));

	mux_2level_tapbuf_size2 mux_left_track_57 (
		.in({chany_top_in[122], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_34_sram_inv[0:1]),
		.out(chanx_left_out[28]));

	mux_2level_tapbuf_size2 mux_left_track_59 (
		.in({chany_top_in[121], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_35_sram_inv[0:1]),
		.out(chanx_left_out[29]));

	mux_2level_tapbuf_size2 mux_left_track_77 (
		.in({chany_top_in[112], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_36_sram_inv[0:1]),
		.out(chanx_left_out[38]));

	mux_2level_tapbuf_size2 mux_left_track_79 (
		.in({chany_top_in[111], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_37_sram_inv[0:1]),
		.out(chanx_left_out[39]));

	mux_2level_tapbuf_size2 mux_left_track_97 (
		.in({chany_top_in[102], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_38_sram_inv[0:1]),
		.out(chanx_left_out[48]));

	mux_2level_tapbuf_size2 mux_left_track_99 (
		.in({chany_top_in[101], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_39_sram_inv[0:1]),
		.out(chanx_left_out[49]));

	mux_2level_tapbuf_size2 mux_left_track_117 (
		.in({chany_top_in[92], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_40_sram_inv[0:1]),
		.out(chanx_left_out[58]));

	mux_2level_tapbuf_size2 mux_left_track_119 (
		.in({chany_top_in[91], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_41_sram_inv[0:1]),
		.out(chanx_left_out[59]));

	mux_2level_tapbuf_size2 mux_left_track_137 (
		.in({chany_top_in[82], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_42_sram_inv[0:1]),
		.out(chanx_left_out[68]));

	mux_2level_tapbuf_size2 mux_left_track_139 (
		.in({chany_top_in[81], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_43_sram_inv[0:1]),
		.out(chanx_left_out[69]));

	mux_2level_tapbuf_size2 mux_left_track_157 (
		.in({chany_top_in[72], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_44_sram_inv[0:1]),
		.out(chanx_left_out[78]));

	mux_2level_tapbuf_size2 mux_left_track_159 (
		.in({chany_top_in[71], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_45_sram_inv[0:1]),
		.out(chanx_left_out[79]));

	mux_2level_tapbuf_size2 mux_left_track_177 (
		.in({chany_top_in[62], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_46_sram_inv[0:1]),
		.out(chanx_left_out[88]));

	mux_2level_tapbuf_size2 mux_left_track_179 (
		.in({chany_top_in[61], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_47_sram_inv[0:1]),
		.out(chanx_left_out[89]));

	mux_2level_tapbuf_size2 mux_left_track_197 (
		.in({chany_top_in[52], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_48_sram_inv[0:1]),
		.out(chanx_left_out[98]));

	mux_2level_tapbuf_size2 mux_left_track_199 (
		.in({chany_top_in[51], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_49_sram_inv[0:1]),
		.out(chanx_left_out[99]));

	mux_2level_tapbuf_size2 mux_left_track_217 (
		.in({chany_top_in[42], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_50_sram_inv[0:1]),
		.out(chanx_left_out[108]));

	mux_2level_tapbuf_size2 mux_left_track_219 (
		.in({chany_top_in[41], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_51_sram_inv[0:1]),
		.out(chanx_left_out[109]));

	mux_2level_tapbuf_size2 mux_left_track_237 (
		.in({chany_top_in[32], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_52_sram_inv[0:1]),
		.out(chanx_left_out[118]));

	mux_2level_tapbuf_size2 mux_left_track_239 (
		.in({chany_top_in[31], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_53_sram_inv[0:1]),
		.out(chanx_left_out[119]));

	mux_2level_tapbuf_size2 mux_left_track_257 (
		.in({chany_top_in[22], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_54_sram_inv[0:1]),
		.out(chanx_left_out[128]));

	mux_2level_tapbuf_size2 mux_left_track_259 (
		.in({chany_top_in[21], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_55_sram_inv[0:1]),
		.out(chanx_left_out[129]));

	mux_2level_tapbuf_size2 mux_left_track_277 (
		.in({chany_top_in[12], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_56_sram_inv[0:1]),
		.out(chanx_left_out[138]));

	mux_2level_tapbuf_size2 mux_left_track_279 (
		.in({chany_top_in[11], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_57_sram_inv[0:1]),
		.out(chanx_left_out[139]));

	mux_2level_tapbuf_size2 mux_left_track_297 (
		.in({chany_top_in[2], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_58_sram_inv[0:1]),
		.out(chanx_left_out[148]));

	mux_2level_tapbuf_size2 mux_left_track_299 (
		.in({chany_top_in[1], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_59_sram_inv[0:1]),
		.out(chanx_left_out[149]));

	mux_2level_tapbuf_size2_mem mem_top_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_0_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_1_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_2_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_38 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_3_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_4_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_5_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_6_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_78 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_7_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_8_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_9_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_10_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_118 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_11_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_12_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_138 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_13_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_14_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_158 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_15_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_16_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_178 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_17_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_196 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_79_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_18_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_198 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_19_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_87_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_20_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_218 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_21_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_236 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_95_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_22_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_238 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_23_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_103_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_24_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_258 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_25_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_276 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_111_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_26_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_278 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_27_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_119_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_28_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_298 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_29_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_127_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_30_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_19 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_31_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_37 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_135_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_32_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_39 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_33_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_143_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_34_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_59 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_35_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_77 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_151_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_36_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_79 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_37_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_97 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_159_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_38_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_99 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_39_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_117 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_167_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_40_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_119 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_41_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_137 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_175_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_42_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_139 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_43_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_157 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_183_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_44_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_159 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_45_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_177 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_191_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_46_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_179 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_47_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_197 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_199_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_48_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_199 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_49_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_217 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_207_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_50_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_219 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_51_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_237 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_215_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_52_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_239 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_53_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_257 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_223_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_54_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_259 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_55_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_277 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_231_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_56_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_279 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_57_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_297 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_239_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_58_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_left_track_299 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_59_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_11__0_ -----

//----- Default net type -----
// `default_nettype wire



