/home/bas33767/Desktop/DD_Lab_exercise/OpenFPGA/Fabric/ihp-sg13g2/libs.ref/sg13g2_stdcell/lef/sg13g2_stdcell.lef