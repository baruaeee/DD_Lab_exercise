//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Mon Jul  7 22:56:04 2025
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for fpga_top -----
module fpga_top(op_clk,
                op_reset,
                op_set,
                pReset,
                prog_clk,
                gfpga_pad_GPIO_PAD,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] op_clk;
//----- GLOBAL PORTS -----
input [0:0] op_reset;
//----- GLOBAL PORTS -----
input [0:0] op_set;
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GPIO PORTS -----
inout [0:223] gfpga_pad_GPIO_PAD;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__undriven_ccff_head;
wire [0:0] cbx_1__0__undriven_ccff_tail;
wire [0:149] cbx_1__0__undriven_chanx_left_in;
wire [0:149] cbx_1__0__undriven_chanx_left_out;
wire [0:149] cbx_1__0__undriven_chanx_right_in;
wire [0:149] cbx_1__0__undriven_chanx_right_out;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_1__1__undriven_ccff_head;
wire [0:0] cbx_1__1__undriven_ccff_tail;
wire [0:149] cbx_1__1__undriven_chanx_left_in;
wire [0:149] cbx_1__1__undriven_chanx_left_out;
wire [0:149] cbx_1__1__undriven_chanx_right_in;
wire [0:149] cbx_1__1__undriven_chanx_right_out;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_1__2__undriven_ccff_head;
wire [0:0] cbx_1__2__undriven_ccff_tail;
wire [0:149] cbx_1__2__undriven_chanx_left_in;
wire [0:149] cbx_1__2__undriven_chanx_left_out;
wire [0:149] cbx_1__2__undriven_chanx_right_in;
wire [0:149] cbx_1__2__undriven_chanx_right_out;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_1__3__undriven_ccff_head;
wire [0:0] cbx_1__3__undriven_ccff_tail;
wire [0:149] cbx_1__3__undriven_chanx_left_in;
wire [0:149] cbx_1__3__undriven_chanx_left_out;
wire [0:149] cbx_1__3__undriven_chanx_right_in;
wire [0:149] cbx_1__3__undriven_chanx_right_out;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_1__4__undriven_ccff_head;
wire [0:0] cbx_1__4__undriven_ccff_tail;
wire [0:149] cbx_1__4__undriven_chanx_left_in;
wire [0:149] cbx_1__4__undriven_chanx_left_out;
wire [0:149] cbx_1__4__undriven_chanx_right_in;
wire [0:149] cbx_1__4__undriven_chanx_right_out;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_1__5__undriven_ccff_head;
wire [0:0] cbx_1__5__undriven_ccff_tail;
wire [0:149] cbx_1__5__undriven_chanx_left_in;
wire [0:149] cbx_1__5__undriven_chanx_left_out;
wire [0:149] cbx_1__5__undriven_chanx_right_in;
wire [0:149] cbx_1__5__undriven_chanx_right_out;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_1__6__undriven_ccff_head;
wire [0:0] cbx_1__6__undriven_ccff_tail;
wire [0:149] cbx_1__6__undriven_chanx_left_in;
wire [0:149] cbx_1__6__undriven_chanx_left_out;
wire [0:149] cbx_1__6__undriven_chanx_right_in;
wire [0:149] cbx_1__6__undriven_chanx_right_out;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_1__7__undriven_ccff_head;
wire [0:0] cbx_1__7__undriven_ccff_tail;
wire [0:149] cbx_1__7__undriven_chanx_left_in;
wire [0:149] cbx_1__7__undriven_chanx_left_out;
wire [0:149] cbx_1__7__undriven_chanx_right_in;
wire [0:149] cbx_1__7__undriven_chanx_right_out;
wire [0:0] cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_2__0__undriven_ccff_head;
wire [0:0] cbx_2__0__undriven_ccff_tail;
wire [0:149] cbx_2__0__undriven_chanx_left_in;
wire [0:149] cbx_2__0__undriven_chanx_left_out;
wire [0:149] cbx_2__0__undriven_chanx_right_in;
wire [0:149] cbx_2__0__undriven_chanx_right_out;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_;
wire [0:0] cbx_2__2__undriven_ccff_head;
wire [0:0] cbx_2__2__undriven_ccff_tail;
wire [0:149] cbx_2__2__undriven_chanx_left_in;
wire [0:149] cbx_2__2__undriven_chanx_left_out;
wire [0:149] cbx_2__2__undriven_chanx_right_in;
wire [0:149] cbx_2__2__undriven_chanx_right_out;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_;
wire [0:0] cbx_2__4__undriven_ccff_head;
wire [0:0] cbx_2__4__undriven_ccff_tail;
wire [0:149] cbx_2__4__undriven_chanx_left_in;
wire [0:149] cbx_2__4__undriven_chanx_left_out;
wire [0:149] cbx_2__4__undriven_chanx_right_in;
wire [0:149] cbx_2__4__undriven_chanx_right_out;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_;
wire [0:149] cbx_2__6__undriven_chanx_left_in;
wire [0:149] cbx_2__6__undriven_chanx_left_out;
wire [0:149] cbx_2__6__undriven_chanx_right_in;
wire [0:149] cbx_2__6__undriven_chanx_right_out;
wire [0:0] cbx_2__7__undriven_ccff_head;
wire [0:0] cbx_2__7__undriven_ccff_tail;
wire [0:149] cbx_2__7__undriven_chanx_left_in;
wire [0:149] cbx_2__7__undriven_chanx_left_out;
wire [0:149] cbx_2__7__undriven_chanx_right_in;
wire [0:149] cbx_2__7__undriven_chanx_right_out;
wire [0:0] cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_3__0__undriven_ccff_head;
wire [0:0] cbx_3__0__undriven_ccff_tail;
wire [0:149] cbx_3__0__undriven_chanx_left_in;
wire [0:149] cbx_3__0__undriven_chanx_left_out;
wire [0:149] cbx_3__0__undriven_chanx_right_in;
wire [0:149] cbx_3__0__undriven_chanx_right_out;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_3__1__undriven_ccff_head;
wire [0:0] cbx_3__1__undriven_ccff_tail;
wire [0:149] cbx_3__1__undriven_chanx_left_in;
wire [0:149] cbx_3__1__undriven_chanx_left_out;
wire [0:149] cbx_3__1__undriven_chanx_right_in;
wire [0:149] cbx_3__1__undriven_chanx_right_out;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_3__2__undriven_ccff_head;
wire [0:0] cbx_3__2__undriven_ccff_tail;
wire [0:149] cbx_3__2__undriven_chanx_left_in;
wire [0:149] cbx_3__2__undriven_chanx_left_out;
wire [0:149] cbx_3__2__undriven_chanx_right_in;
wire [0:149] cbx_3__2__undriven_chanx_right_out;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_3__3__undriven_ccff_head;
wire [0:0] cbx_3__3__undriven_ccff_tail;
wire [0:149] cbx_3__3__undriven_chanx_left_in;
wire [0:149] cbx_3__3__undriven_chanx_left_out;
wire [0:149] cbx_3__3__undriven_chanx_right_in;
wire [0:149] cbx_3__3__undriven_chanx_right_out;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_3__4__undriven_ccff_head;
wire [0:0] cbx_3__4__undriven_ccff_tail;
wire [0:149] cbx_3__4__undriven_chanx_left_in;
wire [0:149] cbx_3__4__undriven_chanx_left_out;
wire [0:149] cbx_3__4__undriven_chanx_right_in;
wire [0:149] cbx_3__4__undriven_chanx_right_out;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_3__5__undriven_ccff_head;
wire [0:0] cbx_3__5__undriven_ccff_tail;
wire [0:149] cbx_3__5__undriven_chanx_left_in;
wire [0:149] cbx_3__5__undriven_chanx_left_out;
wire [0:149] cbx_3__5__undriven_chanx_right_in;
wire [0:149] cbx_3__5__undriven_chanx_right_out;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_3__6__undriven_ccff_head;
wire [0:0] cbx_3__6__undriven_ccff_tail;
wire [0:149] cbx_3__6__undriven_chanx_left_in;
wire [0:149] cbx_3__6__undriven_chanx_left_out;
wire [0:149] cbx_3__6__undriven_chanx_right_in;
wire [0:149] cbx_3__6__undriven_chanx_right_out;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_3__7__undriven_ccff_head;
wire [0:0] cbx_3__7__undriven_ccff_tail;
wire [0:149] cbx_3__7__undriven_chanx_left_in;
wire [0:149] cbx_3__7__undriven_chanx_left_out;
wire [0:149] cbx_3__7__undriven_chanx_right_in;
wire [0:149] cbx_3__7__undriven_chanx_right_out;
wire [0:0] cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_4__0__undriven_ccff_head;
wire [0:0] cbx_4__0__undriven_ccff_tail;
wire [0:149] cbx_4__0__undriven_chanx_left_in;
wire [0:149] cbx_4__0__undriven_chanx_left_out;
wire [0:149] cbx_4__0__undriven_chanx_right_in;
wire [0:149] cbx_4__0__undriven_chanx_right_out;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_4__1__undriven_ccff_head;
wire [0:0] cbx_4__1__undriven_ccff_tail;
wire [0:149] cbx_4__1__undriven_chanx_left_in;
wire [0:149] cbx_4__1__undriven_chanx_left_out;
wire [0:149] cbx_4__1__undriven_chanx_right_in;
wire [0:149] cbx_4__1__undriven_chanx_right_out;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_4__2__undriven_ccff_head;
wire [0:0] cbx_4__2__undriven_ccff_tail;
wire [0:149] cbx_4__2__undriven_chanx_left_in;
wire [0:149] cbx_4__2__undriven_chanx_left_out;
wire [0:149] cbx_4__2__undriven_chanx_right_in;
wire [0:149] cbx_4__2__undriven_chanx_right_out;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_4__3__undriven_ccff_head;
wire [0:0] cbx_4__3__undriven_ccff_tail;
wire [0:149] cbx_4__3__undriven_chanx_left_in;
wire [0:149] cbx_4__3__undriven_chanx_left_out;
wire [0:149] cbx_4__3__undriven_chanx_right_in;
wire [0:149] cbx_4__3__undriven_chanx_right_out;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_4__4__undriven_ccff_head;
wire [0:0] cbx_4__4__undriven_ccff_tail;
wire [0:149] cbx_4__4__undriven_chanx_left_in;
wire [0:149] cbx_4__4__undriven_chanx_left_out;
wire [0:149] cbx_4__4__undriven_chanx_right_in;
wire [0:149] cbx_4__4__undriven_chanx_right_out;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_4__5__undriven_ccff_head;
wire [0:0] cbx_4__5__undriven_ccff_tail;
wire [0:149] cbx_4__5__undriven_chanx_left_in;
wire [0:149] cbx_4__5__undriven_chanx_left_out;
wire [0:149] cbx_4__5__undriven_chanx_right_in;
wire [0:149] cbx_4__5__undriven_chanx_right_out;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_4__6__undriven_ccff_head;
wire [0:0] cbx_4__6__undriven_ccff_tail;
wire [0:149] cbx_4__6__undriven_chanx_left_in;
wire [0:149] cbx_4__6__undriven_chanx_left_out;
wire [0:149] cbx_4__6__undriven_chanx_right_in;
wire [0:149] cbx_4__6__undriven_chanx_right_out;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_4__7__undriven_ccff_head;
wire [0:0] cbx_4__7__undriven_ccff_tail;
wire [0:149] cbx_4__7__undriven_chanx_left_in;
wire [0:149] cbx_4__7__undriven_chanx_left_out;
wire [0:149] cbx_4__7__undriven_chanx_right_in;
wire [0:149] cbx_4__7__undriven_chanx_right_out;
wire [0:0] cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_5__0__undriven_ccff_head;
wire [0:0] cbx_5__0__undriven_ccff_tail;
wire [0:149] cbx_5__0__undriven_chanx_left_in;
wire [0:149] cbx_5__0__undriven_chanx_left_out;
wire [0:149] cbx_5__0__undriven_chanx_right_in;
wire [0:149] cbx_5__0__undriven_chanx_right_out;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_5__1__undriven_ccff_head;
wire [0:0] cbx_5__1__undriven_ccff_tail;
wire [0:149] cbx_5__1__undriven_chanx_left_in;
wire [0:149] cbx_5__1__undriven_chanx_left_out;
wire [0:149] cbx_5__1__undriven_chanx_right_in;
wire [0:149] cbx_5__1__undriven_chanx_right_out;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_5__2__undriven_ccff_head;
wire [0:0] cbx_5__2__undriven_ccff_tail;
wire [0:149] cbx_5__2__undriven_chanx_left_in;
wire [0:149] cbx_5__2__undriven_chanx_left_out;
wire [0:149] cbx_5__2__undriven_chanx_right_in;
wire [0:149] cbx_5__2__undriven_chanx_right_out;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_5__3__undriven_ccff_head;
wire [0:0] cbx_5__3__undriven_ccff_tail;
wire [0:149] cbx_5__3__undriven_chanx_left_in;
wire [0:149] cbx_5__3__undriven_chanx_left_out;
wire [0:149] cbx_5__3__undriven_chanx_right_in;
wire [0:149] cbx_5__3__undriven_chanx_right_out;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_5__4__undriven_ccff_head;
wire [0:0] cbx_5__4__undriven_ccff_tail;
wire [0:149] cbx_5__4__undriven_chanx_left_in;
wire [0:149] cbx_5__4__undriven_chanx_left_out;
wire [0:149] cbx_5__4__undriven_chanx_right_in;
wire [0:149] cbx_5__4__undriven_chanx_right_out;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_5__5__undriven_ccff_head;
wire [0:0] cbx_5__5__undriven_ccff_tail;
wire [0:149] cbx_5__5__undriven_chanx_left_in;
wire [0:149] cbx_5__5__undriven_chanx_left_out;
wire [0:149] cbx_5__5__undriven_chanx_right_in;
wire [0:149] cbx_5__5__undriven_chanx_right_out;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_5__6__undriven_ccff_head;
wire [0:0] cbx_5__6__undriven_ccff_tail;
wire [0:149] cbx_5__6__undriven_chanx_left_in;
wire [0:149] cbx_5__6__undriven_chanx_left_out;
wire [0:149] cbx_5__6__undriven_chanx_right_in;
wire [0:149] cbx_5__6__undriven_chanx_right_out;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_5__7__undriven_ccff_head;
wire [0:0] cbx_5__7__undriven_ccff_tail;
wire [0:149] cbx_5__7__undriven_chanx_left_in;
wire [0:149] cbx_5__7__undriven_chanx_left_out;
wire [0:149] cbx_5__7__undriven_chanx_right_in;
wire [0:149] cbx_5__7__undriven_chanx_right_out;
wire [0:0] cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_6__0__undriven_ccff_head;
wire [0:0] cbx_6__0__undriven_ccff_tail;
wire [0:149] cbx_6__0__undriven_chanx_left_in;
wire [0:149] cbx_6__0__undriven_chanx_left_out;
wire [0:149] cbx_6__0__undriven_chanx_right_in;
wire [0:149] cbx_6__0__undriven_chanx_right_out;
wire [0:0] cbx_6__6__undriven_ccff_head;
wire [0:0] cbx_6__6__undriven_ccff_tail;
wire [0:149] cbx_6__6__undriven_chanx_left_in;
wire [0:149] cbx_6__6__undriven_chanx_left_out;
wire [0:149] cbx_6__6__undriven_chanx_right_in;
wire [0:149] cbx_6__6__undriven_chanx_right_out;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_6__7__undriven_ccff_head;
wire [0:0] cbx_6__7__undriven_ccff_tail;
wire [0:149] cbx_6__7__undriven_chanx_left_in;
wire [0:149] cbx_6__7__undriven_chanx_left_out;
wire [0:149] cbx_6__7__undriven_chanx_right_in;
wire [0:149] cbx_6__7__undriven_chanx_right_out;
wire [0:0] cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_7__0__undriven_ccff_head;
wire [0:0] cbx_7__0__undriven_ccff_tail;
wire [0:149] cbx_7__0__undriven_chanx_left_in;
wire [0:149] cbx_7__0__undriven_chanx_left_out;
wire [0:149] cbx_7__0__undriven_chanx_right_in;
wire [0:149] cbx_7__0__undriven_chanx_right_out;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_7__1__undriven_ccff_head;
wire [0:0] cbx_7__1__undriven_ccff_tail;
wire [0:149] cbx_7__1__undriven_chanx_left_in;
wire [0:149] cbx_7__1__undriven_chanx_left_out;
wire [0:149] cbx_7__1__undriven_chanx_right_in;
wire [0:149] cbx_7__1__undriven_chanx_right_out;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_7__2__undriven_ccff_head;
wire [0:0] cbx_7__2__undriven_ccff_tail;
wire [0:149] cbx_7__2__undriven_chanx_left_in;
wire [0:149] cbx_7__2__undriven_chanx_left_out;
wire [0:149] cbx_7__2__undriven_chanx_right_in;
wire [0:149] cbx_7__2__undriven_chanx_right_out;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_7__3__undriven_ccff_head;
wire [0:0] cbx_7__3__undriven_ccff_tail;
wire [0:149] cbx_7__3__undriven_chanx_left_in;
wire [0:149] cbx_7__3__undriven_chanx_left_out;
wire [0:149] cbx_7__3__undriven_chanx_right_in;
wire [0:149] cbx_7__3__undriven_chanx_right_out;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_7__4__undriven_ccff_head;
wire [0:0] cbx_7__4__undriven_ccff_tail;
wire [0:149] cbx_7__4__undriven_chanx_left_in;
wire [0:149] cbx_7__4__undriven_chanx_left_out;
wire [0:149] cbx_7__4__undriven_chanx_right_in;
wire [0:149] cbx_7__4__undriven_chanx_right_out;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_7__5__undriven_ccff_head;
wire [0:0] cbx_7__5__undriven_ccff_tail;
wire [0:149] cbx_7__5__undriven_chanx_left_in;
wire [0:149] cbx_7__5__undriven_chanx_left_out;
wire [0:149] cbx_7__5__undriven_chanx_right_in;
wire [0:149] cbx_7__5__undriven_chanx_right_out;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_7__6__undriven_ccff_head;
wire [0:0] cbx_7__6__undriven_ccff_tail;
wire [0:149] cbx_7__6__undriven_chanx_left_in;
wire [0:149] cbx_7__6__undriven_chanx_left_out;
wire [0:149] cbx_7__6__undriven_chanx_right_in;
wire [0:149] cbx_7__6__undriven_chanx_right_out;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_7__7__undriven_ccff_head;
wire [0:0] cbx_7__7__undriven_ccff_tail;
wire [0:149] cbx_7__7__undriven_chanx_left_in;
wire [0:149] cbx_7__7__undriven_chanx_left_out;
wire [0:149] cbx_7__7__undriven_chanx_right_in;
wire [0:149] cbx_7__7__undriven_chanx_right_out;
wire [0:0] cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__undriven_ccff_head;
wire [0:0] cby_0__1__undriven_ccff_tail;
wire [0:149] cby_0__1__undriven_chany_bottom_in;
wire [0:149] cby_0__1__undriven_chany_bottom_out;
wire [0:149] cby_0__1__undriven_chany_top_in;
wire [0:149] cby_0__1__undriven_chany_top_out;
wire [0:0] cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__2__undriven_ccff_head;
wire [0:0] cby_0__2__undriven_ccff_tail;
wire [0:149] cby_0__2__undriven_chany_bottom_in;
wire [0:149] cby_0__2__undriven_chany_bottom_out;
wire [0:149] cby_0__2__undriven_chany_top_in;
wire [0:149] cby_0__2__undriven_chany_top_out;
wire [0:0] cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__3__undriven_ccff_head;
wire [0:0] cby_0__3__undriven_ccff_tail;
wire [0:149] cby_0__3__undriven_chany_bottom_in;
wire [0:149] cby_0__3__undriven_chany_bottom_out;
wire [0:149] cby_0__3__undriven_chany_top_in;
wire [0:149] cby_0__3__undriven_chany_top_out;
wire [0:0] cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__4__undriven_ccff_head;
wire [0:0] cby_0__4__undriven_ccff_tail;
wire [0:149] cby_0__4__undriven_chany_bottom_in;
wire [0:149] cby_0__4__undriven_chany_bottom_out;
wire [0:149] cby_0__4__undriven_chany_top_in;
wire [0:149] cby_0__4__undriven_chany_top_out;
wire [0:0] cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__5__undriven_ccff_head;
wire [0:0] cby_0__5__undriven_ccff_tail;
wire [0:149] cby_0__5__undriven_chany_bottom_in;
wire [0:149] cby_0__5__undriven_chany_bottom_out;
wire [0:149] cby_0__5__undriven_chany_top_in;
wire [0:149] cby_0__5__undriven_chany_top_out;
wire [0:0] cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__6__undriven_ccff_head;
wire [0:0] cby_0__6__undriven_ccff_tail;
wire [0:149] cby_0__6__undriven_chany_bottom_in;
wire [0:149] cby_0__6__undriven_chany_bottom_out;
wire [0:149] cby_0__6__undriven_chany_top_in;
wire [0:149] cby_0__6__undriven_chany_top_out;
wire [0:0] cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__7__undriven_ccff_head;
wire [0:0] cby_0__7__undriven_ccff_tail;
wire [0:149] cby_0__7__undriven_chany_bottom_in;
wire [0:149] cby_0__7__undriven_chany_bottom_out;
wire [0:149] cby_0__7__undriven_chany_top_in;
wire [0:149] cby_0__7__undriven_chany_top_out;
wire [0:0] cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_1__1__undriven_ccff_head;
wire [0:0] cby_1__1__undriven_ccff_tail;
wire [0:149] cby_1__1__undriven_chany_bottom_in;
wire [0:149] cby_1__1__undriven_chany_bottom_out;
wire [0:149] cby_1__1__undriven_chany_top_in;
wire [0:149] cby_1__1__undriven_chany_top_out;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__2__undriven_ccff_head;
wire [0:0] cby_1__2__undriven_ccff_tail;
wire [0:149] cby_1__2__undriven_chany_bottom_in;
wire [0:149] cby_1__2__undriven_chany_bottom_out;
wire [0:149] cby_1__2__undriven_chany_top_in;
wire [0:149] cby_1__2__undriven_chany_top_out;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__undriven_ccff_head;
wire [0:0] cby_1__3__undriven_ccff_tail;
wire [0:149] cby_1__3__undriven_chany_bottom_in;
wire [0:149] cby_1__3__undriven_chany_bottom_out;
wire [0:149] cby_1__3__undriven_chany_top_in;
wire [0:149] cby_1__3__undriven_chany_top_out;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__4__undriven_ccff_head;
wire [0:0] cby_1__4__undriven_ccff_tail;
wire [0:149] cby_1__4__undriven_chany_bottom_in;
wire [0:149] cby_1__4__undriven_chany_bottom_out;
wire [0:149] cby_1__4__undriven_chany_top_in;
wire [0:149] cby_1__4__undriven_chany_top_out;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__undriven_ccff_head;
wire [0:0] cby_1__5__undriven_ccff_tail;
wire [0:149] cby_1__5__undriven_chany_bottom_in;
wire [0:149] cby_1__5__undriven_chany_bottom_out;
wire [0:149] cby_1__5__undriven_chany_top_in;
wire [0:149] cby_1__5__undriven_chany_top_out;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__6__undriven_ccff_head;
wire [0:0] cby_1__6__undriven_ccff_tail;
wire [0:149] cby_1__6__undriven_chany_bottom_in;
wire [0:149] cby_1__6__undriven_chany_bottom_out;
wire [0:149] cby_1__6__undriven_chany_top_in;
wire [0:149] cby_1__6__undriven_chany_top_out;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__7__undriven_ccff_head;
wire [0:0] cby_1__7__undriven_ccff_tail;
wire [0:149] cby_1__7__undriven_chany_bottom_in;
wire [0:149] cby_1__7__undriven_chany_bottom_out;
wire [0:149] cby_1__7__undriven_chany_top_in;
wire [0:149] cby_1__7__undriven_chany_top_out;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_2__1__undriven_ccff_head;
wire [0:0] cby_2__1__undriven_ccff_tail;
wire [0:149] cby_2__1__undriven_chany_bottom_in;
wire [0:149] cby_2__1__undriven_chany_bottom_out;
wire [0:149] cby_2__1__undriven_chany_top_in;
wire [0:149] cby_2__1__undriven_chany_top_out;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:149] cby_2__2__undriven_chany_bottom_in;
wire [0:149] cby_2__2__undriven_chany_bottom_out;
wire [0:149] cby_2__2__undriven_chany_top_in;
wire [0:149] cby_2__2__undriven_chany_top_out;
wire [0:0] cby_2__3__undriven_ccff_head;
wire [0:0] cby_2__3__undriven_ccff_tail;
wire [0:149] cby_2__3__undriven_chany_bottom_in;
wire [0:149] cby_2__3__undriven_chany_bottom_out;
wire [0:149] cby_2__3__undriven_chany_top_in;
wire [0:149] cby_2__3__undriven_chany_top_out;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:149] cby_2__4__undriven_chany_bottom_in;
wire [0:149] cby_2__4__undriven_chany_bottom_out;
wire [0:149] cby_2__4__undriven_chany_top_in;
wire [0:149] cby_2__4__undriven_chany_top_out;
wire [0:0] cby_2__5__undriven_ccff_head;
wire [0:0] cby_2__5__undriven_ccff_tail;
wire [0:149] cby_2__5__undriven_chany_bottom_in;
wire [0:149] cby_2__5__undriven_chany_bottom_out;
wire [0:149] cby_2__5__undriven_chany_top_in;
wire [0:149] cby_2__5__undriven_chany_top_out;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:149] cby_2__6__undriven_chany_bottom_in;
wire [0:149] cby_2__6__undriven_chany_bottom_out;
wire [0:149] cby_2__6__undriven_chany_top_in;
wire [0:149] cby_2__6__undriven_chany_top_out;
wire [0:149] cby_2__7__undriven_chany_bottom_in;
wire [0:149] cby_2__7__undriven_chany_bottom_out;
wire [0:149] cby_2__7__undriven_chany_top_in;
wire [0:149] cby_2__7__undriven_chany_top_out;
wire [0:0] cby_3__1__undriven_ccff_head;
wire [0:0] cby_3__1__undriven_ccff_tail;
wire [0:149] cby_3__1__undriven_chany_bottom_in;
wire [0:149] cby_3__1__undriven_chany_bottom_out;
wire [0:149] cby_3__1__undriven_chany_top_in;
wire [0:149] cby_3__1__undriven_chany_top_out;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__undriven_ccff_head;
wire [0:0] cby_3__2__undriven_ccff_tail;
wire [0:149] cby_3__2__undriven_chany_bottom_in;
wire [0:149] cby_3__2__undriven_chany_bottom_out;
wire [0:149] cby_3__2__undriven_chany_top_in;
wire [0:149] cby_3__2__undriven_chany_top_out;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__3__undriven_ccff_head;
wire [0:0] cby_3__3__undriven_ccff_tail;
wire [0:149] cby_3__3__undriven_chany_bottom_in;
wire [0:149] cby_3__3__undriven_chany_bottom_out;
wire [0:149] cby_3__3__undriven_chany_top_in;
wire [0:149] cby_3__3__undriven_chany_top_out;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__4__undriven_ccff_head;
wire [0:0] cby_3__4__undriven_ccff_tail;
wire [0:149] cby_3__4__undriven_chany_bottom_in;
wire [0:149] cby_3__4__undriven_chany_bottom_out;
wire [0:149] cby_3__4__undriven_chany_top_in;
wire [0:149] cby_3__4__undriven_chany_top_out;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__5__undriven_ccff_head;
wire [0:0] cby_3__5__undriven_ccff_tail;
wire [0:149] cby_3__5__undriven_chany_bottom_in;
wire [0:149] cby_3__5__undriven_chany_bottom_out;
wire [0:149] cby_3__5__undriven_chany_top_in;
wire [0:149] cby_3__5__undriven_chany_top_out;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__6__undriven_ccff_head;
wire [0:0] cby_3__6__undriven_ccff_tail;
wire [0:149] cby_3__6__undriven_chany_bottom_in;
wire [0:149] cby_3__6__undriven_chany_bottom_out;
wire [0:149] cby_3__6__undriven_chany_top_in;
wire [0:149] cby_3__6__undriven_chany_top_out;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__7__undriven_ccff_head;
wire [0:0] cby_3__7__undriven_ccff_tail;
wire [0:149] cby_3__7__undriven_chany_bottom_in;
wire [0:149] cby_3__7__undriven_chany_bottom_out;
wire [0:149] cby_3__7__undriven_chany_top_in;
wire [0:149] cby_3__7__undriven_chany_top_out;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_4__1__undriven_ccff_head;
wire [0:0] cby_4__1__undriven_ccff_tail;
wire [0:149] cby_4__1__undriven_chany_bottom_in;
wire [0:149] cby_4__1__undriven_chany_bottom_out;
wire [0:149] cby_4__1__undriven_chany_top_in;
wire [0:149] cby_4__1__undriven_chany_top_out;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_4__2__undriven_ccff_head;
wire [0:0] cby_4__2__undriven_ccff_tail;
wire [0:149] cby_4__2__undriven_chany_bottom_in;
wire [0:149] cby_4__2__undriven_chany_bottom_out;
wire [0:149] cby_4__2__undriven_chany_top_in;
wire [0:149] cby_4__2__undriven_chany_top_out;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_4__3__undriven_ccff_head;
wire [0:0] cby_4__3__undriven_ccff_tail;
wire [0:149] cby_4__3__undriven_chany_bottom_in;
wire [0:149] cby_4__3__undriven_chany_bottom_out;
wire [0:149] cby_4__3__undriven_chany_top_in;
wire [0:149] cby_4__3__undriven_chany_top_out;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_4__4__undriven_ccff_head;
wire [0:0] cby_4__4__undriven_ccff_tail;
wire [0:149] cby_4__4__undriven_chany_bottom_in;
wire [0:149] cby_4__4__undriven_chany_bottom_out;
wire [0:149] cby_4__4__undriven_chany_top_in;
wire [0:149] cby_4__4__undriven_chany_top_out;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_4__5__undriven_ccff_head;
wire [0:0] cby_4__5__undriven_ccff_tail;
wire [0:149] cby_4__5__undriven_chany_bottom_in;
wire [0:149] cby_4__5__undriven_chany_bottom_out;
wire [0:149] cby_4__5__undriven_chany_top_in;
wire [0:149] cby_4__5__undriven_chany_top_out;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_4__6__undriven_ccff_head;
wire [0:0] cby_4__6__undriven_ccff_tail;
wire [0:149] cby_4__6__undriven_chany_bottom_in;
wire [0:149] cby_4__6__undriven_chany_bottom_out;
wire [0:149] cby_4__6__undriven_chany_top_in;
wire [0:149] cby_4__6__undriven_chany_top_out;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_4__7__undriven_ccff_head;
wire [0:0] cby_4__7__undriven_ccff_tail;
wire [0:149] cby_4__7__undriven_chany_bottom_in;
wire [0:149] cby_4__7__undriven_chany_bottom_out;
wire [0:149] cby_4__7__undriven_chany_top_in;
wire [0:149] cby_4__7__undriven_chany_top_out;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_5__1__undriven_ccff_head;
wire [0:0] cby_5__1__undriven_ccff_tail;
wire [0:149] cby_5__1__undriven_chany_bottom_in;
wire [0:149] cby_5__1__undriven_chany_bottom_out;
wire [0:149] cby_5__1__undriven_chany_top_in;
wire [0:149] cby_5__1__undriven_chany_top_out;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_19_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_20_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_21_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_22_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_23_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_24_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_25_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_26_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_27_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_28_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_29_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_30_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_31_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_32_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_33_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_34_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_35_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] cby_5__2__undriven_ccff_head;
wire [0:0] cby_5__2__undriven_ccff_tail;
wire [0:149] cby_5__2__undriven_chany_bottom_in;
wire [0:149] cby_5__2__undriven_chany_bottom_out;
wire [0:149] cby_5__2__undriven_chany_top_in;
wire [0:149] cby_5__2__undriven_chany_top_out;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_5__3__undriven_ccff_head;
wire [0:0] cby_5__3__undriven_ccff_tail;
wire [0:149] cby_5__3__undriven_chany_bottom_in;
wire [0:149] cby_5__3__undriven_chany_bottom_out;
wire [0:149] cby_5__3__undriven_chany_top_in;
wire [0:149] cby_5__3__undriven_chany_top_out;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_5__4__undriven_ccff_head;
wire [0:0] cby_5__4__undriven_ccff_tail;
wire [0:149] cby_5__4__undriven_chany_bottom_in;
wire [0:149] cby_5__4__undriven_chany_bottom_out;
wire [0:149] cby_5__4__undriven_chany_top_in;
wire [0:149] cby_5__4__undriven_chany_top_out;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_5__5__undriven_ccff_head;
wire [0:0] cby_5__5__undriven_ccff_tail;
wire [0:149] cby_5__5__undriven_chany_bottom_in;
wire [0:149] cby_5__5__undriven_chany_bottom_out;
wire [0:149] cby_5__5__undriven_chany_top_in;
wire [0:149] cby_5__5__undriven_chany_top_out;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_5__6__undriven_ccff_head;
wire [0:0] cby_5__6__undriven_ccff_tail;
wire [0:149] cby_5__6__undriven_chany_bottom_in;
wire [0:149] cby_5__6__undriven_chany_bottom_out;
wire [0:149] cby_5__6__undriven_chany_top_in;
wire [0:149] cby_5__6__undriven_chany_top_out;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_5__7__undriven_ccff_head;
wire [0:0] cby_5__7__undriven_ccff_tail;
wire [0:149] cby_5__7__undriven_chany_bottom_in;
wire [0:149] cby_5__7__undriven_chany_bottom_out;
wire [0:149] cby_5__7__undriven_chany_top_in;
wire [0:149] cby_5__7__undriven_chany_top_out;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_6__1__undriven_ccff_head;
wire [0:0] cby_6__1__undriven_ccff_tail;
wire [0:149] cby_6__1__undriven_chany_bottom_in;
wire [0:149] cby_6__1__undriven_chany_bottom_out;
wire [0:149] cby_6__1__undriven_chany_top_in;
wire [0:149] cby_6__1__undriven_chany_top_out;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_19_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_20_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_21_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_22_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_23_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_24_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_25_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_26_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_27_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_28_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_29_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_30_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_31_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_32_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_33_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_34_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_35_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_9_;
wire [0:149] cby_6__2__undriven_chany_bottom_in;
wire [0:149] cby_6__2__undriven_chany_bottom_out;
wire [0:149] cby_6__2__undriven_chany_top_in;
wire [0:149] cby_6__2__undriven_chany_top_out;
wire [0:149] cby_6__3__undriven_chany_bottom_in;
wire [0:149] cby_6__3__undriven_chany_bottom_out;
wire [0:149] cby_6__3__undriven_chany_top_in;
wire [0:149] cby_6__3__undriven_chany_top_out;
wire [0:149] cby_6__4__undriven_chany_bottom_in;
wire [0:149] cby_6__4__undriven_chany_bottom_out;
wire [0:149] cby_6__4__undriven_chany_top_in;
wire [0:149] cby_6__4__undriven_chany_top_out;
wire [0:149] cby_6__5__undriven_chany_bottom_in;
wire [0:149] cby_6__5__undriven_chany_bottom_out;
wire [0:149] cby_6__5__undriven_chany_top_in;
wire [0:149] cby_6__5__undriven_chany_top_out;
wire [0:149] cby_6__6__undriven_chany_bottom_in;
wire [0:149] cby_6__6__undriven_chany_bottom_out;
wire [0:149] cby_6__6__undriven_chany_top_in;
wire [0:149] cby_6__6__undriven_chany_top_out;
wire [0:0] cby_6__7__undriven_ccff_head;
wire [0:0] cby_6__7__undriven_ccff_tail;
wire [0:149] cby_6__7__undriven_chany_bottom_in;
wire [0:149] cby_6__7__undriven_chany_bottom_out;
wire [0:149] cby_6__7__undriven_chany_top_in;
wire [0:149] cby_6__7__undriven_chany_top_out;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_7__1__undriven_ccff_head;
wire [0:0] cby_7__1__undriven_ccff_tail;
wire [0:149] cby_7__1__undriven_chany_bottom_in;
wire [0:149] cby_7__1__undriven_chany_bottom_out;
wire [0:149] cby_7__1__undriven_chany_top_in;
wire [0:149] cby_7__1__undriven_chany_top_out;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_7__2__undriven_ccff_head;
wire [0:0] cby_7__2__undriven_ccff_tail;
wire [0:149] cby_7__2__undriven_chany_bottom_in;
wire [0:149] cby_7__2__undriven_chany_bottom_out;
wire [0:149] cby_7__2__undriven_chany_top_in;
wire [0:149] cby_7__2__undriven_chany_top_out;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_7__3__undriven_ccff_head;
wire [0:0] cby_7__3__undriven_ccff_tail;
wire [0:149] cby_7__3__undriven_chany_bottom_in;
wire [0:149] cby_7__3__undriven_chany_bottom_out;
wire [0:149] cby_7__3__undriven_chany_top_in;
wire [0:149] cby_7__3__undriven_chany_top_out;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_7__4__undriven_ccff_head;
wire [0:0] cby_7__4__undriven_ccff_tail;
wire [0:149] cby_7__4__undriven_chany_bottom_in;
wire [0:149] cby_7__4__undriven_chany_bottom_out;
wire [0:149] cby_7__4__undriven_chany_top_in;
wire [0:149] cby_7__4__undriven_chany_top_out;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_7__5__undriven_ccff_head;
wire [0:0] cby_7__5__undriven_ccff_tail;
wire [0:149] cby_7__5__undriven_chany_bottom_in;
wire [0:149] cby_7__5__undriven_chany_bottom_out;
wire [0:149] cby_7__5__undriven_chany_top_in;
wire [0:149] cby_7__5__undriven_chany_top_out;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_7__6__undriven_ccff_head;
wire [0:0] cby_7__6__undriven_ccff_tail;
wire [0:149] cby_7__6__undriven_chany_bottom_in;
wire [0:149] cby_7__6__undriven_chany_bottom_out;
wire [0:149] cby_7__6__undriven_chany_top_in;
wire [0:149] cby_7__6__undriven_chany_top_out;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_7__7__undriven_ccff_head;
wire [0:0] cby_7__7__undriven_ccff_tail;
wire [0:149] cby_7__7__undriven_chany_bottom_in;
wire [0:149] cby_7__7__undriven_chany_bottom_out;
wire [0:149] cby_7__7__undriven_chany_top_in;
wire [0:149] cby_7__7__undriven_chany_top_out;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_1__1__undriven_ccff_head;
wire [0:0] grid_clb_1__1__undriven_ccff_tail;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_1__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_1__2__undriven_ccff_head;
wire [0:0] grid_clb_1__2__undriven_ccff_tail;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_1__3__undriven_ccff_head;
wire [0:0] grid_clb_1__3__undriven_ccff_tail;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_1__3__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_1__4__undriven_ccff_head;
wire [0:0] grid_clb_1__4__undriven_ccff_tail;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_1__4__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_1__5__undriven_ccff_head;
wire [0:0] grid_clb_1__5__undriven_ccff_tail;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_1__5__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_1__6__undriven_ccff_head;
wire [0:0] grid_clb_1__6__undriven_ccff_tail;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_1__6__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_1__7__undriven_ccff_head;
wire [0:0] grid_clb_1__7__undriven_ccff_tail;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_1__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_3__1__undriven_ccff_head;
wire [0:0] grid_clb_3__1__undriven_ccff_tail;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_3__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_3__2__undriven_ccff_head;
wire [0:0] grid_clb_3__2__undriven_ccff_tail;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_3__3__undriven_ccff_head;
wire [0:0] grid_clb_3__3__undriven_ccff_tail;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_3__3__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_3__4__undriven_ccff_head;
wire [0:0] grid_clb_3__4__undriven_ccff_tail;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_3__4__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_3__5__undriven_ccff_head;
wire [0:0] grid_clb_3__5__undriven_ccff_tail;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_3__5__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_3__6__undriven_ccff_head;
wire [0:0] grid_clb_3__6__undriven_ccff_tail;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_3__6__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_3__7__undriven_ccff_head;
wire [0:0] grid_clb_3__7__undriven_ccff_tail;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_3__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_4__1__undriven_ccff_head;
wire [0:0] grid_clb_4__1__undriven_ccff_tail;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_4__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_4__2__undriven_ccff_head;
wire [0:0] grid_clb_4__2__undriven_ccff_tail;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_4__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_4__3__undriven_ccff_head;
wire [0:0] grid_clb_4__3__undriven_ccff_tail;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_4__3__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_4__4__undriven_ccff_head;
wire [0:0] grid_clb_4__4__undriven_ccff_tail;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_4__4__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_4__5__undriven_ccff_head;
wire [0:0] grid_clb_4__5__undriven_ccff_tail;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_4__5__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_4__6__undriven_ccff_head;
wire [0:0] grid_clb_4__6__undriven_ccff_tail;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_4__6__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_4__7__undriven_ccff_head;
wire [0:0] grid_clb_4__7__undriven_ccff_tail;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_4__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_5__1__undriven_ccff_head;
wire [0:0] grid_clb_5__1__undriven_ccff_tail;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_5__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_5__2__undriven_ccff_head;
wire [0:0] grid_clb_5__2__undriven_ccff_tail;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_5__3__undriven_ccff_head;
wire [0:0] grid_clb_5__3__undriven_ccff_tail;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_5__3__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_5__4__undriven_ccff_head;
wire [0:0] grid_clb_5__4__undriven_ccff_tail;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_5__4__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_5__5__undriven_ccff_head;
wire [0:0] grid_clb_5__5__undriven_ccff_tail;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_5__5__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_5__6__undriven_ccff_head;
wire [0:0] grid_clb_5__6__undriven_ccff_tail;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_5__6__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_5__7__undriven_ccff_head;
wire [0:0] grid_clb_5__7__undriven_ccff_tail;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_5__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_6__7__undriven_ccff_head;
wire [0:0] grid_clb_6__7__undriven_ccff_tail;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_6__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_7__1__undriven_ccff_head;
wire [0:0] grid_clb_7__1__undriven_ccff_tail;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_7__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_7__2__undriven_ccff_head;
wire [0:0] grid_clb_7__2__undriven_ccff_tail;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_7__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_7__3__undriven_ccff_head;
wire [0:0] grid_clb_7__3__undriven_ccff_tail;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_7__3__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_7__4__undriven_ccff_head;
wire [0:0] grid_clb_7__4__undriven_ccff_tail;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_7__4__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_7__5__undriven_ccff_head;
wire [0:0] grid_clb_7__5__undriven_ccff_tail;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_7__5__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_7__6__undriven_ccff_head;
wire [0:0] grid_clb_7__6__undriven_ccff_tail;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_7__6__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_7__7__undriven_ccff_head;
wire [0:0] grid_clb_7__7__undriven_ccff_tail;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_7__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_io_bottom_1__0__undriven_ccff_head;
wire [0:0] grid_io_bottom_1__0__undriven_ccff_tail;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_ccff_head;
wire [0:0] grid_io_bottom_2__0__undriven_ccff_tail;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_ccff_head;
wire [0:0] grid_io_bottom_3__0__undriven_ccff_tail;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_ccff_head;
wire [0:0] grid_io_bottom_4__0__undriven_ccff_tail;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_ccff_head;
wire [0:0] grid_io_bottom_5__0__undriven_ccff_tail;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_ccff_head;
wire [0:0] grid_io_bottom_6__0__undriven_ccff_tail;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_ccff_head;
wire [0:0] grid_io_bottom_7__0__undriven_ccff_tail;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_left_0__1__undriven_ccff_head;
wire [0:0] grid_io_left_0__1__undriven_ccff_tail;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0__1__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_left_0__2__undriven_ccff_head;
wire [0:0] grid_io_left_0__2__undriven_ccff_tail;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0__2__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_left_0__3__undriven_ccff_head;
wire [0:0] grid_io_left_0__3__undriven_ccff_tail;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0__3__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_left_0__4__undriven_ccff_head;
wire [0:0] grid_io_left_0__4__undriven_ccff_tail;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0__4__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_left_0__5__undriven_ccff_head;
wire [0:0] grid_io_left_0__5__undriven_ccff_tail;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0__5__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_left_0__6__undriven_ccff_head;
wire [0:0] grid_io_left_0__6__undriven_ccff_tail;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0__6__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_left_0__7__undriven_ccff_head;
wire [0:0] grid_io_left_0__7__undriven_ccff_tail;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0__7__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_right_8__1__undriven_ccff_head;
wire [0:0] grid_io_right_8__1__undriven_ccff_tail;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_8__1__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_right_8__2__undriven_ccff_head;
wire [0:0] grid_io_right_8__2__undriven_ccff_tail;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_8__2__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_right_8__3__undriven_ccff_head;
wire [0:0] grid_io_right_8__3__undriven_ccff_tail;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_8__3__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_right_8__4__undriven_ccff_head;
wire [0:0] grid_io_right_8__4__undriven_ccff_tail;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_8__4__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_right_8__5__undriven_ccff_head;
wire [0:0] grid_io_right_8__5__undriven_ccff_tail;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_8__5__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_right_8__6__undriven_ccff_head;
wire [0:0] grid_io_right_8__6__undriven_ccff_tail;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_8__6__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_right_8__7__undriven_ccff_head;
wire [0:0] grid_io_right_8__7__undriven_ccff_tail;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_8__7__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_top_1__8__undriven_ccff_head;
wire [0:0] grid_io_top_1__8__undriven_ccff_tail;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_top_2__8__undriven_ccff_head;
wire [0:0] grid_io_top_2__8__undriven_ccff_tail;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_top_3__8__undriven_ccff_head;
wire [0:0] grid_io_top_3__8__undriven_ccff_tail;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_top_4__8__undriven_ccff_head;
wire [0:0] grid_io_top_4__8__undriven_ccff_tail;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_top_5__8__undriven_ccff_head;
wire [0:0] grid_io_top_5__8__undriven_ccff_tail;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_top_6__8__undriven_ccff_head;
wire [0:0] grid_io_top_6__8__undriven_ccff_tail;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_io_top_7__8__undriven_ccff_head;
wire [0:0] grid_io_top_7__8__undriven_ccff_tail;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_5_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_7_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_4_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_5_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_6_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_7_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_6_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_8_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_9_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_ren_0_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_5_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_7_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_9_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_in_1_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_in_3_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_out_0_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_out_1_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_out_2_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_out_3_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_raddr_0_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_raddr_2_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_raddr_4_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_waddr_1_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_waddr_3_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_5_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_7_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_4_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_5_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_6_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_7_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_6_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_8_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_9_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_ren_0_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_5_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_7_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_9_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_in_1_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_in_3_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_out_0_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_out_1_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_out_2_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_out_3_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_raddr_0_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_raddr_2_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_raddr_4_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_waddr_1_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_waddr_3_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_5_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_7_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_4_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_5_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_6_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_7_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_6_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_8_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_9_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_ren_0_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_5_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_7_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_9_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_in_1_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_in_3_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_out_0_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_out_1_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_out_2_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_out_3_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_raddr_0_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_raddr_2_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_raddr_4_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_waddr_1_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_waddr_3_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] grid_mult_36_6__1__undriven_ccff_head;
wire [0:0] grid_mult_36_6__1__undriven_ccff_tail;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_19_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_20_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_21_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_22_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_23_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_24_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_25_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_26_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_27_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_28_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_29_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_30_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_31_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_32_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_33_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_34_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_35_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_38_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_39_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_40_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_41_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_42_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_43_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_44_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_45_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_46_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_47_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_48_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_49_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_50_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_51_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_52_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_53_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_54_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_55_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_56_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_57_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_58_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_59_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_60_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_61_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_62_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_63_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_64_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_65_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_66_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_67_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_68_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_69_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_70_;
wire [0:0] grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_71_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_19_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_20_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_21_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_22_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_23_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_24_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_25_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_26_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_27_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_28_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_29_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_30_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_31_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_32_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_33_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_34_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_35_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_9_;
wire [0:0] sb_0__0__undriven_ccff_head;
wire [0:0] sb_0__0__undriven_ccff_tail;
wire [0:149] sb_0__0__undriven_chanx_right_in;
wire [0:149] sb_0__0__undriven_chanx_right_out;
wire [0:149] sb_0__0__undriven_chany_top_in;
wire [0:149] sb_0__0__undriven_chany_top_out;
wire [0:0] sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_ccff_head;
wire [0:0] sb_0__1__undriven_ccff_tail;
wire [0:149] sb_0__1__undriven_chanx_right_in;
wire [0:149] sb_0__1__undriven_chanx_right_out;
wire [0:149] sb_0__1__undriven_chany_bottom_in;
wire [0:149] sb_0__1__undriven_chany_bottom_out;
wire [0:149] sb_0__1__undriven_chany_top_in;
wire [0:149] sb_0__1__undriven_chany_top_out;
wire [0:0] sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_ccff_head;
wire [0:0] sb_0__2__undriven_ccff_tail;
wire [0:149] sb_0__2__undriven_chanx_right_in;
wire [0:149] sb_0__2__undriven_chanx_right_out;
wire [0:149] sb_0__2__undriven_chany_bottom_in;
wire [0:149] sb_0__2__undriven_chany_bottom_out;
wire [0:149] sb_0__2__undriven_chany_top_in;
wire [0:149] sb_0__2__undriven_chany_top_out;
wire [0:0] sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_ccff_head;
wire [0:0] sb_0__3__undriven_ccff_tail;
wire [0:149] sb_0__3__undriven_chanx_right_in;
wire [0:149] sb_0__3__undriven_chanx_right_out;
wire [0:149] sb_0__3__undriven_chany_bottom_in;
wire [0:149] sb_0__3__undriven_chany_bottom_out;
wire [0:149] sb_0__3__undriven_chany_top_in;
wire [0:149] sb_0__3__undriven_chany_top_out;
wire [0:0] sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_ccff_head;
wire [0:0] sb_0__4__undriven_ccff_tail;
wire [0:149] sb_0__4__undriven_chanx_right_in;
wire [0:149] sb_0__4__undriven_chanx_right_out;
wire [0:149] sb_0__4__undriven_chany_bottom_in;
wire [0:149] sb_0__4__undriven_chany_bottom_out;
wire [0:149] sb_0__4__undriven_chany_top_in;
wire [0:149] sb_0__4__undriven_chany_top_out;
wire [0:0] sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_ccff_head;
wire [0:0] sb_0__5__undriven_ccff_tail;
wire [0:149] sb_0__5__undriven_chanx_right_in;
wire [0:149] sb_0__5__undriven_chanx_right_out;
wire [0:149] sb_0__5__undriven_chany_bottom_in;
wire [0:149] sb_0__5__undriven_chany_bottom_out;
wire [0:149] sb_0__5__undriven_chany_top_in;
wire [0:149] sb_0__5__undriven_chany_top_out;
wire [0:0] sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_ccff_head;
wire [0:0] sb_0__6__undriven_ccff_tail;
wire [0:149] sb_0__6__undriven_chanx_right_in;
wire [0:149] sb_0__6__undriven_chanx_right_out;
wire [0:149] sb_0__6__undriven_chany_bottom_in;
wire [0:149] sb_0__6__undriven_chany_bottom_out;
wire [0:149] sb_0__6__undriven_chany_top_in;
wire [0:149] sb_0__6__undriven_chany_top_out;
wire [0:0] sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_ccff_head;
wire [0:0] sb_0__7__undriven_ccff_tail;
wire [0:149] sb_0__7__undriven_chanx_right_in;
wire [0:149] sb_0__7__undriven_chanx_right_out;
wire [0:149] sb_0__7__undriven_chany_bottom_in;
wire [0:149] sb_0__7__undriven_chany_bottom_out;
wire [0:0] sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_ccff_head;
wire [0:0] sb_1__0__undriven_ccff_tail;
wire [0:149] sb_1__0__undriven_chanx_left_in;
wire [0:149] sb_1__0__undriven_chanx_left_out;
wire [0:149] sb_1__0__undriven_chanx_right_in;
wire [0:149] sb_1__0__undriven_chanx_right_out;
wire [0:149] sb_1__0__undriven_chany_top_in;
wire [0:149] sb_1__0__undriven_chany_top_out;
wire [0:0] sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_1__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_;
wire [0:0] sb_1__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_;
wire [0:0] sb_1__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_;
wire [0:0] sb_1__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_;
wire [0:0] sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__1__undriven_ccff_head;
wire [0:0] sb_1__1__undriven_ccff_tail;
wire [0:149] sb_1__1__undriven_chanx_left_in;
wire [0:149] sb_1__1__undriven_chanx_left_out;
wire [0:149] sb_1__1__undriven_chany_bottom_in;
wire [0:149] sb_1__1__undriven_chany_bottom_out;
wire [0:149] sb_1__1__undriven_chany_top_in;
wire [0:149] sb_1__1__undriven_chany_top_out;
wire [0:0] sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__2__undriven_ccff_head;
wire [0:0] sb_1__2__undriven_ccff_tail;
wire [0:149] sb_1__2__undriven_chanx_left_in;
wire [0:149] sb_1__2__undriven_chanx_left_out;
wire [0:149] sb_1__2__undriven_chanx_right_in;
wire [0:149] sb_1__2__undriven_chanx_right_out;
wire [0:149] sb_1__2__undriven_chany_bottom_in;
wire [0:149] sb_1__2__undriven_chany_bottom_out;
wire [0:149] sb_1__2__undriven_chany_top_in;
wire [0:149] sb_1__2__undriven_chany_top_out;
wire [0:0] sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_1__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_;
wire [0:0] sb_1__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_;
wire [0:0] sb_1__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_;
wire [0:0] sb_1__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_;
wire [0:0] sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__3__undriven_ccff_head;
wire [0:0] sb_1__3__undriven_ccff_tail;
wire [0:149] sb_1__3__undriven_chanx_left_in;
wire [0:149] sb_1__3__undriven_chanx_left_out;
wire [0:149] sb_1__3__undriven_chany_bottom_in;
wire [0:149] sb_1__3__undriven_chany_bottom_out;
wire [0:149] sb_1__3__undriven_chany_top_in;
wire [0:149] sb_1__3__undriven_chany_top_out;
wire [0:0] sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__4__undriven_ccff_head;
wire [0:0] sb_1__4__undriven_ccff_tail;
wire [0:149] sb_1__4__undriven_chanx_left_in;
wire [0:149] sb_1__4__undriven_chanx_left_out;
wire [0:149] sb_1__4__undriven_chanx_right_in;
wire [0:149] sb_1__4__undriven_chanx_right_out;
wire [0:149] sb_1__4__undriven_chany_bottom_in;
wire [0:149] sb_1__4__undriven_chany_bottom_out;
wire [0:149] sb_1__4__undriven_chany_top_in;
wire [0:149] sb_1__4__undriven_chany_top_out;
wire [0:0] sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_1__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_;
wire [0:0] sb_1__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_;
wire [0:0] sb_1__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_;
wire [0:0] sb_1__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_;
wire [0:0] sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__5__undriven_ccff_head;
wire [0:0] sb_1__5__undriven_ccff_tail;
wire [0:149] sb_1__5__undriven_chanx_left_in;
wire [0:149] sb_1__5__undriven_chanx_left_out;
wire [0:149] sb_1__5__undriven_chany_bottom_in;
wire [0:149] sb_1__5__undriven_chany_bottom_out;
wire [0:149] sb_1__5__undriven_chany_top_in;
wire [0:149] sb_1__5__undriven_chany_top_out;
wire [0:0] sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__6__undriven_ccff_head;
wire [0:0] sb_1__6__undriven_ccff_tail;
wire [0:149] sb_1__6__undriven_chanx_left_in;
wire [0:149] sb_1__6__undriven_chanx_left_out;
wire [0:149] sb_1__6__undriven_chanx_right_in;
wire [0:149] sb_1__6__undriven_chanx_right_out;
wire [0:149] sb_1__6__undriven_chany_bottom_in;
wire [0:149] sb_1__6__undriven_chany_bottom_out;
wire [0:149] sb_1__6__undriven_chany_top_in;
wire [0:149] sb_1__6__undriven_chany_top_out;
wire [0:0] sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_1__7__undriven_ccff_head;
wire [0:0] sb_1__7__undriven_ccff_tail;
wire [0:149] sb_1__7__undriven_chanx_left_in;
wire [0:149] sb_1__7__undriven_chanx_left_out;
wire [0:149] sb_1__7__undriven_chanx_right_in;
wire [0:149] sb_1__7__undriven_chanx_right_out;
wire [0:149] sb_1__7__undriven_chany_bottom_in;
wire [0:149] sb_1__7__undriven_chany_bottom_out;
wire [0:0] sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_ccff_head;
wire [0:0] sb_2__0__undriven_ccff_tail;
wire [0:149] sb_2__0__undriven_chanx_left_in;
wire [0:149] sb_2__0__undriven_chanx_left_out;
wire [0:149] sb_2__0__undriven_chanx_right_in;
wire [0:149] sb_2__0__undriven_chanx_right_out;
wire [0:149] sb_2__0__undriven_chany_top_in;
wire [0:149] sb_2__0__undriven_chany_top_out;
wire [0:0] sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_;
wire [0:0] sb_2__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_;
wire [0:0] sb_2__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_;
wire [0:0] sb_2__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_;
wire [0:0] sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_2__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_;
wire [0:0] sb_2__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_;
wire [0:0] sb_2__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_;
wire [0:0] sb_2__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_;
wire [0:0] sb_2__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_;
wire [0:0] sb_2__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_;
wire [0:0] sb_2__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_;
wire [0:0] sb_2__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_;
wire [0:0] sb_2__1__undriven_ccff_head;
wire [0:0] sb_2__1__undriven_ccff_tail;
wire [0:149] sb_2__1__undriven_chanx_right_in;
wire [0:149] sb_2__1__undriven_chanx_right_out;
wire [0:149] sb_2__1__undriven_chany_bottom_in;
wire [0:149] sb_2__1__undriven_chany_bottom_out;
wire [0:149] sb_2__1__undriven_chany_top_in;
wire [0:149] sb_2__1__undriven_chany_top_out;
wire [0:0] sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_2__2__undriven_ccff_head;
wire [0:0] sb_2__2__undriven_ccff_tail;
wire [0:149] sb_2__2__undriven_chanx_left_in;
wire [0:149] sb_2__2__undriven_chanx_left_out;
wire [0:149] sb_2__2__undriven_chanx_right_in;
wire [0:149] sb_2__2__undriven_chanx_right_out;
wire [0:149] sb_2__2__undriven_chany_bottom_in;
wire [0:149] sb_2__2__undriven_chany_bottom_out;
wire [0:149] sb_2__2__undriven_chany_top_in;
wire [0:149] sb_2__2__undriven_chany_top_out;
wire [0:0] sb_2__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_;
wire [0:0] sb_2__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_;
wire [0:0] sb_2__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_;
wire [0:0] sb_2__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_;
wire [0:0] sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_2__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_;
wire [0:0] sb_2__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_;
wire [0:0] sb_2__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_;
wire [0:0] sb_2__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_;
wire [0:0] sb_2__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_;
wire [0:0] sb_2__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_;
wire [0:0] sb_2__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_;
wire [0:0] sb_2__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_;
wire [0:0] sb_2__3__undriven_ccff_head;
wire [0:0] sb_2__3__undriven_ccff_tail;
wire [0:149] sb_2__3__undriven_chanx_right_in;
wire [0:149] sb_2__3__undriven_chanx_right_out;
wire [0:149] sb_2__3__undriven_chany_bottom_in;
wire [0:149] sb_2__3__undriven_chany_bottom_out;
wire [0:149] sb_2__3__undriven_chany_top_in;
wire [0:149] sb_2__3__undriven_chany_top_out;
wire [0:0] sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_2__4__undriven_ccff_head;
wire [0:0] sb_2__4__undriven_ccff_tail;
wire [0:149] sb_2__4__undriven_chanx_left_in;
wire [0:149] sb_2__4__undriven_chanx_left_out;
wire [0:149] sb_2__4__undriven_chanx_right_in;
wire [0:149] sb_2__4__undriven_chanx_right_out;
wire [0:149] sb_2__4__undriven_chany_bottom_in;
wire [0:149] sb_2__4__undriven_chany_bottom_out;
wire [0:149] sb_2__4__undriven_chany_top_in;
wire [0:149] sb_2__4__undriven_chany_top_out;
wire [0:0] sb_2__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_;
wire [0:0] sb_2__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_;
wire [0:0] sb_2__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_;
wire [0:0] sb_2__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_;
wire [0:0] sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_2__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_;
wire [0:0] sb_2__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_;
wire [0:0] sb_2__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_;
wire [0:0] sb_2__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_;
wire [0:0] sb_2__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_;
wire [0:0] sb_2__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_;
wire [0:0] sb_2__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_;
wire [0:0] sb_2__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_;
wire [0:0] sb_2__5__undriven_ccff_head;
wire [0:0] sb_2__5__undriven_ccff_tail;
wire [0:149] sb_2__5__undriven_chanx_right_in;
wire [0:149] sb_2__5__undriven_chanx_right_out;
wire [0:149] sb_2__5__undriven_chany_bottom_in;
wire [0:149] sb_2__5__undriven_chany_bottom_out;
wire [0:149] sb_2__5__undriven_chany_top_in;
wire [0:149] sb_2__5__undriven_chany_top_out;
wire [0:0] sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_2__6__undriven_ccff_head;
wire [0:0] sb_2__6__undriven_ccff_tail;
wire [0:149] sb_2__6__undriven_chanx_left_in;
wire [0:149] sb_2__6__undriven_chanx_left_out;
wire [0:149] sb_2__6__undriven_chanx_right_in;
wire [0:149] sb_2__6__undriven_chanx_right_out;
wire [0:149] sb_2__6__undriven_chany_bottom_in;
wire [0:149] sb_2__6__undriven_chany_bottom_out;
wire [0:149] sb_2__6__undriven_chany_top_in;
wire [0:149] sb_2__6__undriven_chany_top_out;
wire [0:0] sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_2__7__undriven_ccff_head;
wire [0:0] sb_2__7__undriven_ccff_tail;
wire [0:149] sb_2__7__undriven_chanx_left_in;
wire [0:149] sb_2__7__undriven_chanx_left_out;
wire [0:149] sb_2__7__undriven_chanx_right_in;
wire [0:149] sb_2__7__undriven_chanx_right_out;
wire [0:149] sb_2__7__undriven_chany_bottom_in;
wire [0:149] sb_2__7__undriven_chany_bottom_out;
wire [0:0] sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_ccff_head;
wire [0:0] sb_3__0__undriven_ccff_tail;
wire [0:149] sb_3__0__undriven_chanx_left_in;
wire [0:149] sb_3__0__undriven_chanx_left_out;
wire [0:149] sb_3__0__undriven_chanx_right_in;
wire [0:149] sb_3__0__undriven_chanx_right_out;
wire [0:149] sb_3__0__undriven_chany_top_in;
wire [0:149] sb_3__0__undriven_chany_top_out;
wire [0:0] sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__1__undriven_ccff_head;
wire [0:0] sb_3__1__undriven_ccff_tail;
wire [0:149] sb_3__1__undriven_chanx_left_in;
wire [0:149] sb_3__1__undriven_chanx_left_out;
wire [0:149] sb_3__1__undriven_chanx_right_in;
wire [0:149] sb_3__1__undriven_chanx_right_out;
wire [0:149] sb_3__1__undriven_chany_bottom_in;
wire [0:149] sb_3__1__undriven_chany_bottom_out;
wire [0:149] sb_3__1__undriven_chany_top_in;
wire [0:149] sb_3__1__undriven_chany_top_out;
wire [0:0] sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__2__undriven_ccff_head;
wire [0:0] sb_3__2__undriven_ccff_tail;
wire [0:149] sb_3__2__undriven_chanx_left_in;
wire [0:149] sb_3__2__undriven_chanx_left_out;
wire [0:149] sb_3__2__undriven_chanx_right_in;
wire [0:149] sb_3__2__undriven_chanx_right_out;
wire [0:149] sb_3__2__undriven_chany_bottom_in;
wire [0:149] sb_3__2__undriven_chany_bottom_out;
wire [0:149] sb_3__2__undriven_chany_top_in;
wire [0:149] sb_3__2__undriven_chany_top_out;
wire [0:0] sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__3__undriven_ccff_head;
wire [0:0] sb_3__3__undriven_ccff_tail;
wire [0:149] sb_3__3__undriven_chanx_left_in;
wire [0:149] sb_3__3__undriven_chanx_left_out;
wire [0:149] sb_3__3__undriven_chanx_right_in;
wire [0:149] sb_3__3__undriven_chanx_right_out;
wire [0:149] sb_3__3__undriven_chany_bottom_in;
wire [0:149] sb_3__3__undriven_chany_bottom_out;
wire [0:149] sb_3__3__undriven_chany_top_in;
wire [0:149] sb_3__3__undriven_chany_top_out;
wire [0:0] sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__4__undriven_ccff_head;
wire [0:0] sb_3__4__undriven_ccff_tail;
wire [0:149] sb_3__4__undriven_chanx_left_in;
wire [0:149] sb_3__4__undriven_chanx_left_out;
wire [0:149] sb_3__4__undriven_chanx_right_in;
wire [0:149] sb_3__4__undriven_chanx_right_out;
wire [0:149] sb_3__4__undriven_chany_bottom_in;
wire [0:149] sb_3__4__undriven_chany_bottom_out;
wire [0:149] sb_3__4__undriven_chany_top_in;
wire [0:149] sb_3__4__undriven_chany_top_out;
wire [0:0] sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__5__undriven_ccff_head;
wire [0:0] sb_3__5__undriven_ccff_tail;
wire [0:149] sb_3__5__undriven_chanx_left_in;
wire [0:149] sb_3__5__undriven_chanx_left_out;
wire [0:149] sb_3__5__undriven_chanx_right_in;
wire [0:149] sb_3__5__undriven_chanx_right_out;
wire [0:149] sb_3__5__undriven_chany_bottom_in;
wire [0:149] sb_3__5__undriven_chany_bottom_out;
wire [0:149] sb_3__5__undriven_chany_top_in;
wire [0:149] sb_3__5__undriven_chany_top_out;
wire [0:0] sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__6__undriven_ccff_head;
wire [0:0] sb_3__6__undriven_ccff_tail;
wire [0:149] sb_3__6__undriven_chanx_left_in;
wire [0:149] sb_3__6__undriven_chanx_left_out;
wire [0:149] sb_3__6__undriven_chanx_right_in;
wire [0:149] sb_3__6__undriven_chanx_right_out;
wire [0:149] sb_3__6__undriven_chany_bottom_in;
wire [0:149] sb_3__6__undriven_chany_bottom_out;
wire [0:149] sb_3__6__undriven_chany_top_in;
wire [0:149] sb_3__6__undriven_chany_top_out;
wire [0:0] sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_3__7__undriven_ccff_head;
wire [0:0] sb_3__7__undriven_ccff_tail;
wire [0:149] sb_3__7__undriven_chanx_left_in;
wire [0:149] sb_3__7__undriven_chanx_left_out;
wire [0:149] sb_3__7__undriven_chanx_right_in;
wire [0:149] sb_3__7__undriven_chanx_right_out;
wire [0:149] sb_3__7__undriven_chany_bottom_in;
wire [0:149] sb_3__7__undriven_chany_bottom_out;
wire [0:0] sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_ccff_head;
wire [0:0] sb_4__0__undriven_ccff_tail;
wire [0:149] sb_4__0__undriven_chanx_left_in;
wire [0:149] sb_4__0__undriven_chanx_left_out;
wire [0:149] sb_4__0__undriven_chanx_right_in;
wire [0:149] sb_4__0__undriven_chanx_right_out;
wire [0:149] sb_4__0__undriven_chany_top_in;
wire [0:149] sb_4__0__undriven_chany_top_out;
wire [0:0] sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__1__undriven_ccff_head;
wire [0:0] sb_4__1__undriven_ccff_tail;
wire [0:149] sb_4__1__undriven_chanx_left_in;
wire [0:149] sb_4__1__undriven_chanx_left_out;
wire [0:149] sb_4__1__undriven_chanx_right_in;
wire [0:149] sb_4__1__undriven_chanx_right_out;
wire [0:149] sb_4__1__undriven_chany_bottom_in;
wire [0:149] sb_4__1__undriven_chany_bottom_out;
wire [0:149] sb_4__1__undriven_chany_top_in;
wire [0:149] sb_4__1__undriven_chany_top_out;
wire [0:0] sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__2__undriven_ccff_head;
wire [0:0] sb_4__2__undriven_ccff_tail;
wire [0:149] sb_4__2__undriven_chanx_left_in;
wire [0:149] sb_4__2__undriven_chanx_left_out;
wire [0:149] sb_4__2__undriven_chanx_right_in;
wire [0:149] sb_4__2__undriven_chanx_right_out;
wire [0:149] sb_4__2__undriven_chany_bottom_in;
wire [0:149] sb_4__2__undriven_chany_bottom_out;
wire [0:149] sb_4__2__undriven_chany_top_in;
wire [0:149] sb_4__2__undriven_chany_top_out;
wire [0:0] sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__3__undriven_ccff_head;
wire [0:0] sb_4__3__undriven_ccff_tail;
wire [0:149] sb_4__3__undriven_chanx_left_in;
wire [0:149] sb_4__3__undriven_chanx_left_out;
wire [0:149] sb_4__3__undriven_chanx_right_in;
wire [0:149] sb_4__3__undriven_chanx_right_out;
wire [0:149] sb_4__3__undriven_chany_bottom_in;
wire [0:149] sb_4__3__undriven_chany_bottom_out;
wire [0:149] sb_4__3__undriven_chany_top_in;
wire [0:149] sb_4__3__undriven_chany_top_out;
wire [0:0] sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__4__undriven_ccff_head;
wire [0:0] sb_4__4__undriven_ccff_tail;
wire [0:149] sb_4__4__undriven_chanx_left_in;
wire [0:149] sb_4__4__undriven_chanx_left_out;
wire [0:149] sb_4__4__undriven_chanx_right_in;
wire [0:149] sb_4__4__undriven_chanx_right_out;
wire [0:149] sb_4__4__undriven_chany_bottom_in;
wire [0:149] sb_4__4__undriven_chany_bottom_out;
wire [0:149] sb_4__4__undriven_chany_top_in;
wire [0:149] sb_4__4__undriven_chany_top_out;
wire [0:0] sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__5__undriven_ccff_head;
wire [0:0] sb_4__5__undriven_ccff_tail;
wire [0:149] sb_4__5__undriven_chanx_left_in;
wire [0:149] sb_4__5__undriven_chanx_left_out;
wire [0:149] sb_4__5__undriven_chanx_right_in;
wire [0:149] sb_4__5__undriven_chanx_right_out;
wire [0:149] sb_4__5__undriven_chany_bottom_in;
wire [0:149] sb_4__5__undriven_chany_bottom_out;
wire [0:149] sb_4__5__undriven_chany_top_in;
wire [0:149] sb_4__5__undriven_chany_top_out;
wire [0:0] sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__6__undriven_ccff_head;
wire [0:0] sb_4__6__undriven_ccff_tail;
wire [0:149] sb_4__6__undriven_chanx_left_in;
wire [0:149] sb_4__6__undriven_chanx_left_out;
wire [0:149] sb_4__6__undriven_chanx_right_in;
wire [0:149] sb_4__6__undriven_chanx_right_out;
wire [0:149] sb_4__6__undriven_chany_bottom_in;
wire [0:149] sb_4__6__undriven_chany_bottom_out;
wire [0:149] sb_4__6__undriven_chany_top_in;
wire [0:149] sb_4__6__undriven_chany_top_out;
wire [0:0] sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_4__7__undriven_ccff_head;
wire [0:0] sb_4__7__undriven_ccff_tail;
wire [0:149] sb_4__7__undriven_chanx_left_in;
wire [0:149] sb_4__7__undriven_chanx_left_out;
wire [0:149] sb_4__7__undriven_chanx_right_in;
wire [0:149] sb_4__7__undriven_chanx_right_out;
wire [0:149] sb_4__7__undriven_chany_bottom_in;
wire [0:149] sb_4__7__undriven_chany_bottom_out;
wire [0:0] sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_ccff_head;
wire [0:0] sb_5__0__undriven_ccff_tail;
wire [0:149] sb_5__0__undriven_chanx_left_in;
wire [0:149] sb_5__0__undriven_chanx_left_out;
wire [0:149] sb_5__0__undriven_chanx_right_in;
wire [0:149] sb_5__0__undriven_chanx_right_out;
wire [0:149] sb_5__0__undriven_chany_top_in;
wire [0:149] sb_5__0__undriven_chany_top_out;
wire [0:0] sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_38_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_39_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_40_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_41_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_42_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_43_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_44_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_45_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_46_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_47_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_48_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_49_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_50_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_51_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_52_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_53_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_54_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_55_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_56_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_57_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_58_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_59_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_60_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_61_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_62_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_63_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_64_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_65_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_66_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_67_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_68_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_69_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_70_;
wire [0:0] sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_71_;
wire [0:0] sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_38_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_39_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_40_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_41_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_42_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_43_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_44_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_45_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_46_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_47_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_48_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_49_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_50_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_51_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_52_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_53_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_54_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_55_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_56_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_57_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_58_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_59_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_60_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_61_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_62_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_63_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_64_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_65_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_66_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_67_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_68_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_69_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_70_;
wire [0:0] sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_71_;
wire [0:0] sb_5__1__undriven_ccff_head;
wire [0:0] sb_5__1__undriven_ccff_tail;
wire [0:149] sb_5__1__undriven_chanx_left_in;
wire [0:149] sb_5__1__undriven_chanx_left_out;
wire [0:149] sb_5__1__undriven_chany_bottom_in;
wire [0:149] sb_5__1__undriven_chany_bottom_out;
wire [0:149] sb_5__1__undriven_chany_top_in;
wire [0:149] sb_5__1__undriven_chany_top_out;
wire [0:0] sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__2__undriven_ccff_head;
wire [0:0] sb_5__2__undriven_ccff_tail;
wire [0:149] sb_5__2__undriven_chanx_left_in;
wire [0:149] sb_5__2__undriven_chanx_left_out;
wire [0:149] sb_5__2__undriven_chany_bottom_in;
wire [0:149] sb_5__2__undriven_chany_bottom_out;
wire [0:149] sb_5__2__undriven_chany_top_in;
wire [0:149] sb_5__2__undriven_chany_top_out;
wire [0:0] sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__3__undriven_ccff_head;
wire [0:0] sb_5__3__undriven_ccff_tail;
wire [0:149] sb_5__3__undriven_chanx_left_in;
wire [0:149] sb_5__3__undriven_chanx_left_out;
wire [0:149] sb_5__3__undriven_chany_bottom_in;
wire [0:149] sb_5__3__undriven_chany_bottom_out;
wire [0:149] sb_5__3__undriven_chany_top_in;
wire [0:149] sb_5__3__undriven_chany_top_out;
wire [0:0] sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__4__undriven_ccff_head;
wire [0:0] sb_5__4__undriven_ccff_tail;
wire [0:149] sb_5__4__undriven_chanx_left_in;
wire [0:149] sb_5__4__undriven_chanx_left_out;
wire [0:149] sb_5__4__undriven_chany_bottom_in;
wire [0:149] sb_5__4__undriven_chany_bottom_out;
wire [0:149] sb_5__4__undriven_chany_top_in;
wire [0:149] sb_5__4__undriven_chany_top_out;
wire [0:0] sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__5__undriven_ccff_head;
wire [0:0] sb_5__5__undriven_ccff_tail;
wire [0:149] sb_5__5__undriven_chanx_left_in;
wire [0:149] sb_5__5__undriven_chanx_left_out;
wire [0:149] sb_5__5__undriven_chany_bottom_in;
wire [0:149] sb_5__5__undriven_chany_bottom_out;
wire [0:149] sb_5__5__undriven_chany_top_in;
wire [0:149] sb_5__5__undriven_chany_top_out;
wire [0:0] sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__6__undriven_ccff_head;
wire [0:0] sb_5__6__undriven_ccff_tail;
wire [0:149] sb_5__6__undriven_chanx_left_in;
wire [0:149] sb_5__6__undriven_chanx_left_out;
wire [0:149] sb_5__6__undriven_chanx_right_in;
wire [0:149] sb_5__6__undriven_chanx_right_out;
wire [0:149] sb_5__6__undriven_chany_bottom_in;
wire [0:149] sb_5__6__undriven_chany_bottom_out;
wire [0:149] sb_5__6__undriven_chany_top_in;
wire [0:149] sb_5__6__undriven_chany_top_out;
wire [0:0] sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_5__7__undriven_ccff_head;
wire [0:0] sb_5__7__undriven_ccff_tail;
wire [0:149] sb_5__7__undriven_chanx_left_in;
wire [0:149] sb_5__7__undriven_chanx_left_out;
wire [0:149] sb_5__7__undriven_chanx_right_in;
wire [0:149] sb_5__7__undriven_chanx_right_out;
wire [0:149] sb_5__7__undriven_chany_bottom_in;
wire [0:149] sb_5__7__undriven_chany_bottom_out;
wire [0:0] sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_ccff_head;
wire [0:0] sb_6__0__undriven_ccff_tail;
wire [0:149] sb_6__0__undriven_chanx_left_in;
wire [0:149] sb_6__0__undriven_chanx_left_out;
wire [0:149] sb_6__0__undriven_chanx_right_in;
wire [0:149] sb_6__0__undriven_chanx_right_out;
wire [0:149] sb_6__0__undriven_chany_top_in;
wire [0:149] sb_6__0__undriven_chany_top_out;
wire [0:0] sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_9_;
wire [0:0] sb_6__1__undriven_ccff_head;
wire [0:0] sb_6__1__undriven_ccff_tail;
wire [0:149] sb_6__1__undriven_chanx_right_in;
wire [0:149] sb_6__1__undriven_chanx_right_out;
wire [0:149] sb_6__1__undriven_chany_bottom_in;
wire [0:149] sb_6__1__undriven_chany_bottom_out;
wire [0:149] sb_6__1__undriven_chany_top_in;
wire [0:149] sb_6__1__undriven_chany_top_out;
wire [0:0] sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_6__2__undriven_ccff_head;
wire [0:0] sb_6__2__undriven_ccff_tail;
wire [0:149] sb_6__2__undriven_chanx_right_in;
wire [0:149] sb_6__2__undriven_chanx_right_out;
wire [0:149] sb_6__2__undriven_chany_bottom_in;
wire [0:149] sb_6__2__undriven_chany_bottom_out;
wire [0:149] sb_6__2__undriven_chany_top_in;
wire [0:149] sb_6__2__undriven_chany_top_out;
wire [0:0] sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_6__3__undriven_ccff_head;
wire [0:0] sb_6__3__undriven_ccff_tail;
wire [0:149] sb_6__3__undriven_chanx_right_in;
wire [0:149] sb_6__3__undriven_chanx_right_out;
wire [0:149] sb_6__3__undriven_chany_bottom_in;
wire [0:149] sb_6__3__undriven_chany_bottom_out;
wire [0:149] sb_6__3__undriven_chany_top_in;
wire [0:149] sb_6__3__undriven_chany_top_out;
wire [0:0] sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_6__4__undriven_ccff_head;
wire [0:0] sb_6__4__undriven_ccff_tail;
wire [0:149] sb_6__4__undriven_chanx_right_in;
wire [0:149] sb_6__4__undriven_chanx_right_out;
wire [0:149] sb_6__4__undriven_chany_bottom_in;
wire [0:149] sb_6__4__undriven_chany_bottom_out;
wire [0:149] sb_6__4__undriven_chany_top_in;
wire [0:149] sb_6__4__undriven_chany_top_out;
wire [0:0] sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_6__5__undriven_ccff_head;
wire [0:0] sb_6__5__undriven_ccff_tail;
wire [0:149] sb_6__5__undriven_chanx_right_in;
wire [0:149] sb_6__5__undriven_chanx_right_out;
wire [0:149] sb_6__5__undriven_chany_bottom_in;
wire [0:149] sb_6__5__undriven_chany_bottom_out;
wire [0:149] sb_6__5__undriven_chany_top_in;
wire [0:149] sb_6__5__undriven_chany_top_out;
wire [0:0] sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_6__6__undriven_ccff_head;
wire [0:0] sb_6__6__undriven_ccff_tail;
wire [0:149] sb_6__6__undriven_chanx_left_in;
wire [0:149] sb_6__6__undriven_chanx_left_out;
wire [0:149] sb_6__6__undriven_chanx_right_in;
wire [0:149] sb_6__6__undriven_chanx_right_out;
wire [0:149] sb_6__6__undriven_chany_bottom_in;
wire [0:149] sb_6__6__undriven_chany_bottom_out;
wire [0:149] sb_6__6__undriven_chany_top_in;
wire [0:149] sb_6__6__undriven_chany_top_out;
wire [0:0] sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_6__7__undriven_ccff_head;
wire [0:0] sb_6__7__undriven_ccff_tail;
wire [0:149] sb_6__7__undriven_chanx_left_in;
wire [0:149] sb_6__7__undriven_chanx_left_out;
wire [0:149] sb_6__7__undriven_chanx_right_in;
wire [0:149] sb_6__7__undriven_chanx_right_out;
wire [0:149] sb_6__7__undriven_chany_bottom_in;
wire [0:149] sb_6__7__undriven_chany_bottom_out;
wire [0:0] sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_ccff_head;
wire [0:0] sb_7__0__undriven_ccff_tail;
wire [0:149] sb_7__0__undriven_chanx_left_in;
wire [0:149] sb_7__0__undriven_chanx_left_out;
wire [0:149] sb_7__0__undriven_chany_top_in;
wire [0:149] sb_7__0__undriven_chany_top_out;
wire [0:0] sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_ccff_head;
wire [0:0] sb_7__1__undriven_ccff_tail;
wire [0:149] sb_7__1__undriven_chanx_left_in;
wire [0:149] sb_7__1__undriven_chanx_left_out;
wire [0:149] sb_7__1__undriven_chany_bottom_in;
wire [0:149] sb_7__1__undriven_chany_bottom_out;
wire [0:149] sb_7__1__undriven_chany_top_in;
wire [0:149] sb_7__1__undriven_chany_top_out;
wire [0:0] sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_ccff_head;
wire [0:0] sb_7__2__undriven_ccff_tail;
wire [0:149] sb_7__2__undriven_chanx_left_in;
wire [0:149] sb_7__2__undriven_chanx_left_out;
wire [0:149] sb_7__2__undriven_chany_bottom_in;
wire [0:149] sb_7__2__undriven_chany_bottom_out;
wire [0:149] sb_7__2__undriven_chany_top_in;
wire [0:149] sb_7__2__undriven_chany_top_out;
wire [0:0] sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_ccff_head;
wire [0:0] sb_7__3__undriven_ccff_tail;
wire [0:149] sb_7__3__undriven_chanx_left_in;
wire [0:149] sb_7__3__undriven_chanx_left_out;
wire [0:149] sb_7__3__undriven_chany_bottom_in;
wire [0:149] sb_7__3__undriven_chany_bottom_out;
wire [0:149] sb_7__3__undriven_chany_top_in;
wire [0:149] sb_7__3__undriven_chany_top_out;
wire [0:0] sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_ccff_head;
wire [0:0] sb_7__4__undriven_ccff_tail;
wire [0:149] sb_7__4__undriven_chanx_left_in;
wire [0:149] sb_7__4__undriven_chanx_left_out;
wire [0:149] sb_7__4__undriven_chany_bottom_in;
wire [0:149] sb_7__4__undriven_chany_bottom_out;
wire [0:149] sb_7__4__undriven_chany_top_in;
wire [0:149] sb_7__4__undriven_chany_top_out;
wire [0:0] sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_ccff_head;
wire [0:0] sb_7__5__undriven_ccff_tail;
wire [0:149] sb_7__5__undriven_chanx_left_in;
wire [0:149] sb_7__5__undriven_chanx_left_out;
wire [0:149] sb_7__5__undriven_chany_bottom_in;
wire [0:149] sb_7__5__undriven_chany_bottom_out;
wire [0:149] sb_7__5__undriven_chany_top_in;
wire [0:149] sb_7__5__undriven_chany_top_out;
wire [0:0] sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_ccff_head;
wire [0:0] sb_7__6__undriven_ccff_tail;
wire [0:149] sb_7__6__undriven_chanx_left_in;
wire [0:149] sb_7__6__undriven_chanx_left_out;
wire [0:149] sb_7__6__undriven_chany_bottom_in;
wire [0:149] sb_7__6__undriven_chany_bottom_out;
wire [0:149] sb_7__6__undriven_chany_top_in;
wire [0:149] sb_7__6__undriven_chany_top_out;
wire [0:0] sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_ccff_head;
wire [0:0] sb_7__7__undriven_ccff_tail;
wire [0:149] sb_7__7__undriven_chanx_left_in;
wire [0:149] sb_7__7__undriven_chanx_left_out;
wire [0:149] sb_7__7__undriven_chany_bottom_in;
wire [0:149] sb_7__7__undriven_chany_bottom_out;
wire [0:0] sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_io_top grid_io_top_1__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:7]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_1__8__undriven_ccff_head),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_1__8__undriven_ccff_tail));

	grid_io_top grid_io_top_2__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8:15]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_2__8__undriven_ccff_head),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_2__8__undriven_ccff_tail));

	grid_io_top grid_io_top_3__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[16:23]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_3__8__undriven_ccff_head),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_3__8__undriven_ccff_tail));

	grid_io_top grid_io_top_4__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[24:31]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_4__8__undriven_ccff_head),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_4__8__undriven_ccff_tail));

	grid_io_top grid_io_top_5__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[32:39]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_5__8__undriven_ccff_head),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_5__8__undriven_ccff_tail));

	grid_io_top grid_io_top_6__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[40:47]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_6__8__undriven_ccff_head),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_6__8__undriven_ccff_tail));

	grid_io_top grid_io_top_7__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[48:55]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_7__8__undriven_ccff_head),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_7__8__undriven_ccff_tail));

	grid_io_right grid_io_right_8__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[56:63]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_8__7__undriven_ccff_head),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8__7__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_8__7__undriven_ccff_tail));

	grid_io_right grid_io_right_8__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[64:71]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_8__6__undriven_ccff_head),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8__6__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_8__6__undriven_ccff_tail));

	grid_io_right grid_io_right_8__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[72:79]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_8__5__undriven_ccff_head),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8__5__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_8__5__undriven_ccff_tail));

	grid_io_right grid_io_right_8__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[80:87]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_8__4__undriven_ccff_head),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8__4__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_8__4__undriven_ccff_tail));

	grid_io_right grid_io_right_8__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[88:95]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_8__3__undriven_ccff_head),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8__3__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_8__3__undriven_ccff_tail));

	grid_io_right grid_io_right_8__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[96:103]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_8__2__undriven_ccff_head),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8__2__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_8__2__undriven_ccff_tail));

	grid_io_right grid_io_right_8__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[104:111]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_8__1__undriven_ccff_head),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8__1__undriven_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_8__1__undriven_ccff_tail));

	grid_io_bottom grid_io_bottom_7__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[112:119]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_7__0__undriven_ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_7__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_7__0__undriven_ccff_tail));

	grid_io_bottom grid_io_bottom_6__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[120:127]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_6__0__undriven_ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_6__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_6__0__undriven_ccff_tail));

	grid_io_bottom grid_io_bottom_5__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[128:135]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_5__0__undriven_ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_5__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_5__0__undriven_ccff_tail));

	grid_io_bottom grid_io_bottom_4__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[136:143]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_4__0__undriven_ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_4__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_4__0__undriven_ccff_tail));

	grid_io_bottom grid_io_bottom_3__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[144:151]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_3__0__undriven_ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_3__0__undriven_ccff_tail));

	grid_io_bottom grid_io_bottom_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[152:159]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_2__0__undriven_ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_2__0__undriven_ccff_tail));

	grid_io_bottom grid_io_bottom_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[160:167]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_1__0__undriven_ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1__0__undriven_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_1__0__undriven_ccff_tail));

	grid_io_left grid_io_left_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[168:175]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_left_0__1__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0__1__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0__1__undriven_ccff_tail));

	grid_io_left grid_io_left_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[176:183]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_left_0__2__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0__2__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0__2__undriven_ccff_tail));

	grid_io_left grid_io_left_0__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[184:191]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_left_0__3__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0__3__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0__3__undriven_ccff_tail));

	grid_io_left grid_io_left_0__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[192:199]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_left_0__4__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0__4__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0__4__undriven_ccff_tail));

	grid_io_left grid_io_left_0__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[200:207]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_left_0__5__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0__5__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0__5__undriven_ccff_tail));

	grid_io_left grid_io_left_0__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[208:215]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_left_0__6__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0__6__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0__6__undriven_ccff_tail));

	grid_io_left grid_io_left_0__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[216:223]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_left_0__7__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0__7__undriven_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0__7__undriven_ccff_tail));

	grid_clb grid_clb_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_1__1__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1__1__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_1__1__undriven_ccff_tail));

	grid_clb grid_clb_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_1__2__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1__2__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_1__2__undriven_ccff_tail));

	grid_clb grid_clb_1__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__3__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_1__3__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1__3__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_1__3__undriven_ccff_tail));

	grid_clb grid_clb_1__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__4__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_1__4__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1__4__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_1__4__undriven_ccff_tail));

	grid_clb grid_clb_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__5__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_1__5__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1__5__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_1__5__undriven_ccff_tail));

	grid_clb grid_clb_1__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__6__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_1__6__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1__6__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_1__6__undriven_ccff_tail));

	grid_clb grid_clb_1__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_1__7__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_1__7__undriven_ccff_tail));

	grid_clb grid_clb_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_3__1__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3__1__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_3__1__undriven_ccff_tail));

	grid_clb grid_clb_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_3__2__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3__2__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_3__2__undriven_ccff_tail));

	grid_clb grid_clb_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__3__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_3__3__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3__3__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_3__3__undriven_ccff_tail));

	grid_clb grid_clb_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__4__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_3__4__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3__4__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_3__4__undriven_ccff_tail));

	grid_clb grid_clb_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__5__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_3__5__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3__5__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_3__5__undriven_ccff_tail));

	grid_clb grid_clb_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__6__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_3__6__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3__6__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_3__6__undriven_ccff_tail));

	grid_clb grid_clb_3__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_3__7__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_3__7__undriven_ccff_tail));

	grid_clb grid_clb_4__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_4__1__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4__1__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_4__1__undriven_ccff_tail));

	grid_clb grid_clb_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_4__2__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4__2__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_4__2__undriven_ccff_tail));

	grid_clb grid_clb_4__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__3__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_4__3__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4__3__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_4__3__undriven_ccff_tail));

	grid_clb grid_clb_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__4__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_4__4__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4__4__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_4__4__undriven_ccff_tail));

	grid_clb grid_clb_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__5__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_4__5__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4__5__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_4__5__undriven_ccff_tail));

	grid_clb grid_clb_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__6__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_4__6__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4__6__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_4__6__undriven_ccff_tail));

	grid_clb grid_clb_4__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_4__7__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_4__7__undriven_ccff_tail));

	grid_clb grid_clb_5__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_5__1__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5__1__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_5__1__undriven_ccff_tail));

	grid_clb grid_clb_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_5__2__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5__2__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_5__2__undriven_ccff_tail));

	grid_clb grid_clb_5__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__3__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_5__3__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5__3__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_5__3__undriven_ccff_tail));

	grid_clb grid_clb_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__4__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_5__4__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5__4__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_5__4__undriven_ccff_tail));

	grid_clb grid_clb_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__5__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_5__5__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5__5__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_5__5__undriven_ccff_tail));

	grid_clb grid_clb_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__6__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_5__6__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5__6__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_5__6__undriven_ccff_tail));

	grid_clb grid_clb_5__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_5__7__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_5__7__undriven_ccff_tail));

	grid_clb grid_clb_6__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_6__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_6__7__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_6__7__undriven_ccff_tail));

	grid_clb grid_clb_7__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_7__1__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7__1__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_7__1__undriven_ccff_tail));

	grid_clb grid_clb_7__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_7__2__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7__2__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_7__2__undriven_ccff_tail));

	grid_clb grid_clb_7__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__3__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_7__3__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7__3__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_7__3__undriven_ccff_tail));

	grid_clb grid_clb_7__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__4__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_7__4__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7__4__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_7__4__undriven_ccff_tail));

	grid_clb grid_clb_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__5__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_7__5__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7__5__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_7__5__undriven_ccff_tail));

	grid_clb grid_clb_7__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__6__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_7__6__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7__6__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_7__6__undriven_ccff_tail));

	grid_clb grid_clb_7__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_set_0_(op_set),
		.left_width_0_height_0_subtile_0__pin_reset_0_(op_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.ccff_head(grid_clb_7__7__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7__7__undriven_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_7__7__undriven_ccff_tail));

	grid_memory grid_memory_2__1_ (
		.right_width_0_height_0_subtile_0__pin_waddr_0_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_waddr_0_),
		.right_width_0_height_0_subtile_0__pin_waddr_1_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_waddr_1_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_waddr_3_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_waddr_3_),
		.right_width_0_height_0_subtile_0__pin_waddr_4_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_waddr_4_),
		.right_width_0_height_0_subtile_0__pin_raddr_0_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_raddr_0_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_raddr_2_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_raddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_3_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_raddr_3_),
		.right_width_0_height_0_subtile_0__pin_raddr_4_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_raddr_4_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_data_in_1_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_in_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_2_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_in_2_),
		.right_width_0_height_0_subtile_0__pin_data_in_3_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_in_3_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_5_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_6_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_6_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_7_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_7_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_8_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_9_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_9_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_5_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_5_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_6_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_6_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_7_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_8_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_8_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_9_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_9_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_4_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_4_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_5_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_5_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_6_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_6_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_7_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_7_),
		.bottom_width_0_height_0_subtile_0__pin_ren_0_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_ren_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.right_width_0_height_0_subtile_0__pin_data_out_0_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.right_width_0_height_0_subtile_0__pin_data_out_1_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.right_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.right_width_0_height_0_subtile_0__pin_data_out_3_(grid_memory_2__1__undriven_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_5_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_7_(grid_memory_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_7_));

	grid_memory grid_memory_2__3_ (
		.right_width_0_height_0_subtile_0__pin_waddr_0_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_waddr_0_),
		.right_width_0_height_0_subtile_0__pin_waddr_1_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_waddr_1_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_waddr_3_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_waddr_3_),
		.right_width_0_height_0_subtile_0__pin_waddr_4_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_waddr_4_),
		.right_width_0_height_0_subtile_0__pin_raddr_0_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_raddr_0_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_raddr_2_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_raddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_3_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_raddr_3_),
		.right_width_0_height_0_subtile_0__pin_raddr_4_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_raddr_4_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_data_in_1_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_in_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_2_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_in_2_),
		.right_width_0_height_0_subtile_0__pin_data_in_3_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_in_3_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_5_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_6_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_6_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_7_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_7_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_8_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_9_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_9_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_5_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_5_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_6_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_6_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_7_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_8_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_8_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_9_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_9_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_4_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_4_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_5_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_5_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_6_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_6_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_7_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_7_),
		.bottom_width_0_height_0_subtile_0__pin_ren_0_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_ren_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.right_width_0_height_0_subtile_0__pin_data_out_0_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.right_width_0_height_0_subtile_0__pin_data_out_1_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.right_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.right_width_0_height_0_subtile_0__pin_data_out_3_(grid_memory_2__3__undriven_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_5_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_7_(grid_memory_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_7_));

	grid_memory grid_memory_2__5_ (
		.right_width_0_height_0_subtile_0__pin_waddr_0_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_waddr_0_),
		.right_width_0_height_0_subtile_0__pin_waddr_1_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_waddr_1_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_waddr_3_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_waddr_3_),
		.right_width_0_height_0_subtile_0__pin_waddr_4_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_waddr_4_),
		.right_width_0_height_0_subtile_0__pin_raddr_0_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_raddr_0_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_raddr_2_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_raddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_3_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_raddr_3_),
		.right_width_0_height_0_subtile_0__pin_raddr_4_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_raddr_4_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_data_in_1_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_in_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_2_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_in_2_),
		.right_width_0_height_0_subtile_0__pin_data_in_3_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_in_3_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_5_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_6_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_6_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_7_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_7_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_8_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_9_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_waddr_9_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_5_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_5_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_6_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_6_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_7_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_8_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_8_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_9_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_raddr_9_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_4_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_4_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_5_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_5_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_6_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_6_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_7_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_in_7_),
		.bottom_width_0_height_0_subtile_0__pin_ren_0_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_ren_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(op_clk),
		.right_width_0_height_0_subtile_0__pin_data_out_0_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.right_width_0_height_0_subtile_0__pin_data_out_1_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.right_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.right_width_0_height_0_subtile_0__pin_data_out_3_(grid_memory_2__5__undriven_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_5_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_7_(grid_memory_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_data_out_7_));

	grid_mult_36 grid_mult_36_6__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.right_width_0_height_0_subtile_0__pin_a_0_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_0_),
		.right_width_0_height_0_subtile_0__pin_a_1_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_1_),
		.right_width_0_height_0_subtile_0__pin_a_2_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_2_),
		.right_width_0_height_0_subtile_0__pin_a_3_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_3_),
		.right_width_0_height_0_subtile_0__pin_a_4_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_4_),
		.right_width_0_height_0_subtile_0__pin_a_5_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_5_),
		.right_width_0_height_0_subtile_0__pin_a_6_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_6_),
		.right_width_0_height_0_subtile_0__pin_a_7_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_7_),
		.right_width_0_height_0_subtile_0__pin_a_8_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_8_),
		.right_width_0_height_0_subtile_0__pin_a_9_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_9_),
		.right_width_0_height_0_subtile_0__pin_a_10_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_10_),
		.right_width_0_height_0_subtile_0__pin_a_11_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_11_),
		.right_width_0_height_0_subtile_0__pin_a_12_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_12_),
		.right_width_0_height_0_subtile_0__pin_a_13_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_13_),
		.right_width_0_height_0_subtile_0__pin_a_14_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_14_),
		.right_width_0_height_0_subtile_0__pin_a_15_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_15_),
		.right_width_0_height_0_subtile_0__pin_a_16_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_16_),
		.right_width_0_height_0_subtile_0__pin_a_17_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_17_),
		.right_width_0_height_0_subtile_0__pin_a_18_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_18_),
		.right_width_0_height_0_subtile_0__pin_a_19_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_19_),
		.right_width_0_height_0_subtile_0__pin_a_20_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_20_),
		.right_width_0_height_0_subtile_0__pin_a_21_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_21_),
		.right_width_0_height_0_subtile_0__pin_a_22_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_22_),
		.right_width_0_height_0_subtile_0__pin_a_23_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_23_),
		.right_width_0_height_0_subtile_0__pin_a_24_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_24_),
		.right_width_0_height_0_subtile_0__pin_a_25_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_25_),
		.right_width_0_height_0_subtile_0__pin_a_26_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_26_),
		.right_width_0_height_0_subtile_0__pin_a_27_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_27_),
		.right_width_0_height_0_subtile_0__pin_a_28_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_28_),
		.right_width_0_height_0_subtile_0__pin_a_29_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_29_),
		.right_width_0_height_0_subtile_0__pin_a_30_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_30_),
		.right_width_0_height_0_subtile_0__pin_a_31_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_31_),
		.right_width_0_height_0_subtile_0__pin_a_32_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_32_),
		.right_width_0_height_0_subtile_0__pin_a_33_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_33_),
		.right_width_0_height_0_subtile_0__pin_a_34_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_34_),
		.right_width_0_height_0_subtile_0__pin_a_35_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_a_35_),
		.left_width_0_height_0_subtile_0__pin_b_0_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_0_),
		.left_width_0_height_0_subtile_0__pin_b_1_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_1_),
		.left_width_0_height_0_subtile_0__pin_b_2_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_2_),
		.left_width_0_height_0_subtile_0__pin_b_3_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_3_),
		.left_width_0_height_0_subtile_0__pin_b_4_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_4_),
		.left_width_0_height_0_subtile_0__pin_b_5_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_5_),
		.left_width_0_height_0_subtile_0__pin_b_6_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_6_),
		.left_width_0_height_0_subtile_0__pin_b_7_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_7_),
		.left_width_0_height_0_subtile_0__pin_b_8_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_8_),
		.left_width_0_height_0_subtile_0__pin_b_9_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_9_),
		.left_width_0_height_0_subtile_0__pin_b_10_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_10_),
		.left_width_0_height_0_subtile_0__pin_b_11_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_11_),
		.left_width_0_height_0_subtile_0__pin_b_12_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_12_),
		.left_width_0_height_0_subtile_0__pin_b_13_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_13_),
		.left_width_0_height_0_subtile_0__pin_b_14_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_14_),
		.left_width_0_height_0_subtile_0__pin_b_15_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_15_),
		.left_width_0_height_0_subtile_0__pin_b_16_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_16_),
		.left_width_0_height_0_subtile_0__pin_b_17_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_17_),
		.left_width_0_height_0_subtile_0__pin_b_18_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_18_),
		.left_width_0_height_0_subtile_0__pin_b_19_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_19_),
		.left_width_0_height_0_subtile_0__pin_b_20_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_20_),
		.left_width_0_height_0_subtile_0__pin_b_21_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_21_),
		.left_width_0_height_0_subtile_0__pin_b_22_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_22_),
		.left_width_0_height_0_subtile_0__pin_b_23_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_23_),
		.left_width_0_height_0_subtile_0__pin_b_24_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_24_),
		.left_width_0_height_0_subtile_0__pin_b_25_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_25_),
		.left_width_0_height_0_subtile_0__pin_b_26_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_26_),
		.left_width_0_height_0_subtile_0__pin_b_27_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_27_),
		.left_width_0_height_0_subtile_0__pin_b_28_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_28_),
		.left_width_0_height_0_subtile_0__pin_b_29_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_29_),
		.left_width_0_height_0_subtile_0__pin_b_30_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_30_),
		.left_width_0_height_0_subtile_0__pin_b_31_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_31_),
		.left_width_0_height_0_subtile_0__pin_b_32_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_32_),
		.left_width_0_height_0_subtile_0__pin_b_33_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_33_),
		.left_width_0_height_0_subtile_0__pin_b_34_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_34_),
		.left_width_0_height_0_subtile_0__pin_b_35_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_b_35_),
		.ccff_head(grid_mult_36_6__1__undriven_ccff_head),
		.right_width_0_height_0_subtile_0__pin_out_0_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_0_),
		.right_width_0_height_0_subtile_0__pin_out_1_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_1_),
		.right_width_0_height_0_subtile_0__pin_out_2_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_2_),
		.right_width_0_height_0_subtile_0__pin_out_3_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_3_),
		.right_width_0_height_0_subtile_0__pin_out_4_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_4_),
		.right_width_0_height_0_subtile_0__pin_out_5_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_5_),
		.right_width_0_height_0_subtile_0__pin_out_6_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_6_),
		.right_width_0_height_0_subtile_0__pin_out_7_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_7_),
		.right_width_0_height_0_subtile_0__pin_out_8_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_8_),
		.right_width_0_height_0_subtile_0__pin_out_9_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_9_),
		.right_width_0_height_0_subtile_0__pin_out_10_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_10_),
		.right_width_0_height_0_subtile_0__pin_out_11_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_11_),
		.right_width_0_height_0_subtile_0__pin_out_12_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_12_),
		.right_width_0_height_0_subtile_0__pin_out_13_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_13_),
		.right_width_0_height_0_subtile_0__pin_out_14_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_14_),
		.right_width_0_height_0_subtile_0__pin_out_15_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_15_),
		.right_width_0_height_0_subtile_0__pin_out_16_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_16_),
		.right_width_0_height_0_subtile_0__pin_out_17_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_17_),
		.right_width_0_height_0_subtile_0__pin_out_18_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_18_),
		.right_width_0_height_0_subtile_0__pin_out_19_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_19_),
		.right_width_0_height_0_subtile_0__pin_out_20_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_20_),
		.right_width_0_height_0_subtile_0__pin_out_21_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_21_),
		.right_width_0_height_0_subtile_0__pin_out_22_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_22_),
		.right_width_0_height_0_subtile_0__pin_out_23_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_23_),
		.right_width_0_height_0_subtile_0__pin_out_24_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_24_),
		.right_width_0_height_0_subtile_0__pin_out_25_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_25_),
		.right_width_0_height_0_subtile_0__pin_out_26_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_26_),
		.right_width_0_height_0_subtile_0__pin_out_27_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_27_),
		.right_width_0_height_0_subtile_0__pin_out_28_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_28_),
		.right_width_0_height_0_subtile_0__pin_out_29_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_29_),
		.right_width_0_height_0_subtile_0__pin_out_30_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_30_),
		.right_width_0_height_0_subtile_0__pin_out_31_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_31_),
		.right_width_0_height_0_subtile_0__pin_out_32_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_32_),
		.right_width_0_height_0_subtile_0__pin_out_33_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_33_),
		.right_width_0_height_0_subtile_0__pin_out_34_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_34_),
		.right_width_0_height_0_subtile_0__pin_out_35_(grid_mult_36_6__1__undriven_right_width_0_height_0_subtile_0__pin_out_35_),
		.left_width_0_height_0_subtile_0__pin_out_36_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_36_),
		.left_width_0_height_0_subtile_0__pin_out_37_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_37_),
		.left_width_0_height_0_subtile_0__pin_out_38_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_38_),
		.left_width_0_height_0_subtile_0__pin_out_39_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_39_),
		.left_width_0_height_0_subtile_0__pin_out_40_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_40_),
		.left_width_0_height_0_subtile_0__pin_out_41_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_41_),
		.left_width_0_height_0_subtile_0__pin_out_42_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_42_),
		.left_width_0_height_0_subtile_0__pin_out_43_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_43_),
		.left_width_0_height_0_subtile_0__pin_out_44_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_44_),
		.left_width_0_height_0_subtile_0__pin_out_45_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_45_),
		.left_width_0_height_0_subtile_0__pin_out_46_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_46_),
		.left_width_0_height_0_subtile_0__pin_out_47_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_47_),
		.left_width_0_height_0_subtile_0__pin_out_48_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_48_),
		.left_width_0_height_0_subtile_0__pin_out_49_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_49_),
		.left_width_0_height_0_subtile_0__pin_out_50_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_50_),
		.left_width_0_height_0_subtile_0__pin_out_51_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_51_),
		.left_width_0_height_0_subtile_0__pin_out_52_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_52_),
		.left_width_0_height_0_subtile_0__pin_out_53_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_53_),
		.left_width_0_height_0_subtile_0__pin_out_54_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_54_),
		.left_width_0_height_0_subtile_0__pin_out_55_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_55_),
		.left_width_0_height_0_subtile_0__pin_out_56_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_56_),
		.left_width_0_height_0_subtile_0__pin_out_57_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_57_),
		.left_width_0_height_0_subtile_0__pin_out_58_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_58_),
		.left_width_0_height_0_subtile_0__pin_out_59_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_59_),
		.left_width_0_height_0_subtile_0__pin_out_60_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_60_),
		.left_width_0_height_0_subtile_0__pin_out_61_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_61_),
		.left_width_0_height_0_subtile_0__pin_out_62_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_62_),
		.left_width_0_height_0_subtile_0__pin_out_63_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_63_),
		.left_width_0_height_0_subtile_0__pin_out_64_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_64_),
		.left_width_0_height_0_subtile_0__pin_out_65_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_65_),
		.left_width_0_height_0_subtile_0__pin_out_66_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_66_),
		.left_width_0_height_0_subtile_0__pin_out_67_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_67_),
		.left_width_0_height_0_subtile_0__pin_out_68_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_68_),
		.left_width_0_height_0_subtile_0__pin_out_69_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_69_),
		.left_width_0_height_0_subtile_0__pin_out_70_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_70_),
		.left_width_0_height_0_subtile_0__pin_out_71_(grid_mult_36_6__1__undriven_left_width_0_height_0_subtile_0__pin_out_71_),
		.ccff_tail(grid_mult_36_6__1__undriven_ccff_tail));

	sb_0__0_ sb_0__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_0__0__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__0__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(sb_0__0__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_0__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__0__undriven_ccff_head),
		.chany_top_out(sb_0__0__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_0__0__undriven_chanx_right_out[0:149]),
		.ccff_tail(sb_0__0__undriven_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_0__1__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__1__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(sb_0__1__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_0__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_0__1__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__1__undriven_ccff_head),
		.chany_top_out(sb_0__1__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_0__1__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_0__1__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_0__1__undriven_ccff_tail));

	sb_0__1_ sb_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_0__2__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__2__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(sb_0__2__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_0__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_0__2__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__2__undriven_ccff_head),
		.chany_top_out(sb_0__2__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_0__2__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_0__2__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_0__2__undriven_ccff_tail));

	sb_0__1_ sb_0__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_0__3__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__3__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(sb_0__3__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_0__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_0__3__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__3__undriven_ccff_head),
		.chany_top_out(sb_0__3__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_0__3__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_0__3__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_0__3__undriven_ccff_tail));

	sb_0__1_ sb_0__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_0__4__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__4__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(sb_0__4__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_0__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_0__4__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__4__undriven_ccff_head),
		.chany_top_out(sb_0__4__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_0__4__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_0__4__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_0__4__undriven_ccff_tail));

	sb_0__1_ sb_0__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_0__5__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__5__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(sb_0__5__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_0__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_0__5__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__5__undriven_ccff_head),
		.chany_top_out(sb_0__5__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_0__5__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_0__5__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_0__5__undriven_ccff_tail));

	sb_0__1_ sb_0__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_0__6__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__6__undriven_top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(sb_0__6__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_0__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_0__6__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__6__undriven_ccff_head),
		.chany_top_out(sb_0__6__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_0__6__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_0__6__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_0__6__undriven_ccff_tail));

	sb_0__7_ sb_0__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(sb_0__7__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_0__7__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(sb_0__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__7__undriven_ccff_head),
		.chanx_right_out(sb_0__7__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_0__7__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_0__7__undriven_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_1__0__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_1__0__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_(sb_1__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_(sb_1__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_(sb_1__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_(sb_1__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_1__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(sb_1__0__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_1__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_1__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_1__0__undriven_ccff_head),
		.chany_top_out(sb_1__0__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_1__0__undriven_chanx_right_out[0:149]),
		.chanx_left_out(sb_1__0__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_1__0__undriven_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_1__1__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(sb_1__1__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_1__1__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_1__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_1__1__undriven_ccff_head),
		.chany_top_out(sb_1__1__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_1__1__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_1__1__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_1__1__undriven_ccff_tail));

	sb_1__1_ sb_1__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_1__3__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(sb_1__3__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_1__3__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_1__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_1__3__undriven_ccff_head),
		.chany_top_out(sb_1__3__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_1__3__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_1__3__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_1__3__undriven_ccff_tail));

	sb_1__1_ sb_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_1__5__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(sb_1__5__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_1__5__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_1__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_1__5__undriven_ccff_head),
		.chany_top_out(sb_1__5__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_1__5__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_1__5__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_1__5__undriven_ccff_tail));

	sb_1__1_ sb_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_5__2__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(sb_5__2__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_5__2__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_5__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_5__2__undriven_ccff_head),
		.chany_top_out(sb_5__2__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_5__2__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_5__2__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_5__2__undriven_ccff_tail));

	sb_1__1_ sb_5__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_5__3__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(sb_5__3__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_5__3__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_5__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_5__3__undriven_ccff_head),
		.chany_top_out(sb_5__3__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_5__3__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_5__3__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_5__3__undriven_ccff_tail));

	sb_1__1_ sb_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_5__4__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(sb_5__4__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_5__4__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_5__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_5__4__undriven_ccff_head),
		.chany_top_out(sb_5__4__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_5__4__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_5__4__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_5__4__undriven_ccff_tail));

	sb_1__1_ sb_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_5__5__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(sb_5__5__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_5__5__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_5__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_5__5__undriven_ccff_head),
		.chany_top_out(sb_5__5__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_5__5__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_5__5__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_5__5__undriven_ccff_tail));

	sb_1__2_ sb_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_1__2__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_1__2__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_(sb_1__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_(sb_1__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_(sb_1__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_(sb_1__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_),
		.chany_bottom_in(sb_1__2__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_1__2__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_1__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_1__2__undriven_ccff_head),
		.chany_top_out(sb_1__2__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_1__2__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_1__2__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_1__2__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_1__2__undriven_ccff_tail));

	sb_1__2_ sb_1__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_1__4__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_1__4__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_(sb_1__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_(sb_1__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_(sb_1__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_(sb_1__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_),
		.chany_bottom_in(sb_1__4__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_1__4__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_1__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_1__4__undriven_ccff_head),
		.chany_top_out(sb_1__4__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_1__4__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_1__4__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_1__4__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_1__4__undriven_ccff_tail));

	sb_1__6_ sb_1__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_1__6__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_1__6__undriven_chanx_right_in[0:149]),
		.chany_bottom_in(sb_1__6__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_1__6__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_1__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_1__6__undriven_ccff_head),
		.chany_top_out(sb_1__6__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_1__6__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_1__6__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_1__6__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_1__6__undriven_ccff_tail));

	sb_1__7_ sb_1__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(sb_1__7__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_1__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_1__7__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_1__7__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_1__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_1__7__undriven_ccff_head),
		.chanx_right_out(sb_1__7__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_1__7__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_1__7__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_1__7__undriven_ccff_tail));

	sb_1__7_ sb_3__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(sb_3__7__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_3__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_3__7__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_3__7__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_3__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_3__7__undriven_ccff_head),
		.chanx_right_out(sb_3__7__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_3__7__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_3__7__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_3__7__undriven_ccff_tail));

	sb_1__7_ sb_4__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(sb_4__7__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_4__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_4__7__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_4__7__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_4__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_4__7__undriven_ccff_head),
		.chanx_right_out(sb_4__7__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_4__7__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_4__7__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_4__7__undriven_ccff_tail));

	sb_1__7_ sb_5__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(sb_5__7__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_5__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_5__7__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_5__7__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_5__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_5__7__undriven_ccff_head),
		.chanx_right_out(sb_5__7__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_5__7__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_5__7__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_5__7__undriven_ccff_tail));

	sb_1__7_ sb_6__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(sb_6__7__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_6__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_6__7__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_6__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_6__7__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_6__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_6__7__undriven_ccff_head),
		.chanx_right_out(sb_6__7__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_6__7__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_6__7__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_6__7__undriven_ccff_tail));

	sb_2__0_ sb_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_2__0__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_(sb_2__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_(sb_2__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_(sb_2__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_(sb_2__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.chanx_right_in(sb_2__0__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_2__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_2__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(sb_2__0__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_(sb_2__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_(sb_2__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_(sb_2__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_(sb_2__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_2__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_2__0__undriven_ccff_head),
		.chany_top_out(sb_2__0__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_2__0__undriven_chanx_right_out[0:149]),
		.chanx_left_out(sb_2__0__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_2__0__undriven_ccff_tail));

	sb_2__1_ sb_2__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_2__1__undriven_chany_top_in[0:149]),
		.chanx_right_in(sb_2__1__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_2__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_2__1__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_(sb_2__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_(sb_2__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_(sb_2__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_(sb_2__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.ccff_head(sb_2__1__undriven_ccff_head),
		.chany_top_out(sb_2__1__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_2__1__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_2__1__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_2__1__undriven_ccff_tail));

	sb_2__1_ sb_2__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_2__3__undriven_chany_top_in[0:149]),
		.chanx_right_in(sb_2__3__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_2__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_2__3__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_(sb_2__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_(sb_2__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_(sb_2__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_(sb_2__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.ccff_head(sb_2__3__undriven_ccff_head),
		.chany_top_out(sb_2__3__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_2__3__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_2__3__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_2__3__undriven_ccff_tail));

	sb_2__1_ sb_2__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_2__5__undriven_chany_top_in[0:149]),
		.chanx_right_in(sb_2__5__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_2__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_2__5__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_(sb_2__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_(sb_2__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_(sb_2__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_(sb_2__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.ccff_head(sb_2__5__undriven_ccff_head),
		.chany_top_out(sb_2__5__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_2__5__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_2__5__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_2__5__undriven_ccff_tail));

	sb_2__2_ sb_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_2__2__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_(sb_2__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_(sb_2__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_(sb_2__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_(sb_2__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.chanx_right_in(sb_2__2__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_2__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_2__2__undriven_chany_bottom_in[0:149]),
		.chanx_left_in(sb_2__2__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_(sb_2__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_(sb_2__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_(sb_2__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_(sb_2__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_),
		.ccff_head(sb_2__2__undriven_ccff_head),
		.chany_top_out(sb_2__2__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_2__2__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_2__2__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_2__2__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_2__2__undriven_ccff_tail));

	sb_2__2_ sb_2__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_2__4__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_(sb_2__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_(sb_2__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_(sb_2__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_(sb_2__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.chanx_right_in(sb_2__4__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_2__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_2__4__undriven_chany_bottom_in[0:149]),
		.chanx_left_in(sb_2__4__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_(sb_2__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_(sb_2__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_(sb_2__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_(sb_2__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_),
		.ccff_head(sb_2__4__undriven_ccff_head),
		.chany_top_out(sb_2__4__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_2__4__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_2__4__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_2__4__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_2__4__undriven_ccff_tail));

	sb_2__6_ sb_2__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_2__6__undriven_chany_top_in[0:149]),
		.chanx_right_in(sb_2__6__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_2__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_2__6__undriven_chany_bottom_in[0:149]),
		.chanx_left_in(sb_2__6__undriven_chanx_left_in[0:149]),
		.ccff_head(sb_2__6__undriven_ccff_head),
		.chany_top_out(sb_2__6__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_2__6__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_2__6__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_2__6__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_2__6__undriven_ccff_tail));

	sb_2__7_ sb_2__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(sb_2__7__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_2__7__undriven_right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_2__7__undriven_chany_bottom_in[0:149]),
		.chanx_left_in(sb_2__7__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_2__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_2__7__undriven_ccff_head),
		.chanx_right_out(sb_2__7__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_2__7__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_2__7__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_2__7__undriven_ccff_tail));

	sb_3__0_ sb_3__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_3__0__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_3__0__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_3__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(sb_3__0__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_3__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_3__0__undriven_ccff_head),
		.chany_top_out(sb_3__0__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_3__0__undriven_chanx_right_out[0:149]),
		.chanx_left_out(sb_3__0__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_3__0__undriven_ccff_tail));

	sb_3__0_ sb_4__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_4__0__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_4__0__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_4__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(sb_4__0__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_4__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_4__0__undriven_ccff_head),
		.chany_top_out(sb_4__0__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_4__0__undriven_chanx_right_out[0:149]),
		.chanx_left_out(sb_4__0__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_4__0__undriven_ccff_tail));

	sb_3__1_ sb_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_3__1__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_3__1__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_3__1__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_3__1__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_3__1__undriven_ccff_head),
		.chany_top_out(sb_3__1__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_3__1__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_3__1__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_3__1__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_3__1__undriven_ccff_tail));

	sb_3__1_ sb_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_3__2__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_3__2__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_3__2__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_3__2__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_3__2__undriven_ccff_head),
		.chany_top_out(sb_3__2__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_3__2__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_3__2__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_3__2__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_3__2__undriven_ccff_tail));

	sb_3__1_ sb_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_3__3__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_3__3__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_3__3__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_3__3__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_3__3__undriven_ccff_head),
		.chany_top_out(sb_3__3__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_3__3__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_3__3__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_3__3__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_3__3__undriven_ccff_tail));

	sb_3__1_ sb_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_3__4__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_3__4__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_3__4__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_3__4__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_3__4__undriven_ccff_head),
		.chany_top_out(sb_3__4__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_3__4__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_3__4__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_3__4__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_3__4__undriven_ccff_tail));

	sb_3__1_ sb_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_3__5__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_3__5__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_3__5__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_3__5__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_3__5__undriven_ccff_head),
		.chany_top_out(sb_3__5__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_3__5__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_3__5__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_3__5__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_3__5__undriven_ccff_tail));

	sb_3__1_ sb_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_3__6__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_3__6__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_3__6__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_3__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_3__6__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_3__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_3__6__undriven_ccff_head),
		.chany_top_out(sb_3__6__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_3__6__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_3__6__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_3__6__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_3__6__undriven_ccff_tail));

	sb_3__1_ sb_4__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_4__1__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_4__1__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_4__1__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_4__1__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_4__1__undriven_ccff_head),
		.chany_top_out(sb_4__1__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_4__1__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_4__1__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_4__1__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_4__1__undriven_ccff_tail));

	sb_3__1_ sb_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_4__2__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_4__2__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_4__2__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_4__2__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_4__2__undriven_ccff_head),
		.chany_top_out(sb_4__2__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_4__2__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_4__2__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_4__2__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_4__2__undriven_ccff_tail));

	sb_3__1_ sb_4__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_4__3__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_4__3__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_4__3__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_4__3__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_4__3__undriven_ccff_head),
		.chany_top_out(sb_4__3__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_4__3__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_4__3__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_4__3__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_4__3__undriven_ccff_tail));

	sb_3__1_ sb_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_4__4__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_4__4__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_4__4__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_4__4__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_4__4__undriven_ccff_head),
		.chany_top_out(sb_4__4__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_4__4__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_4__4__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_4__4__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_4__4__undriven_ccff_tail));

	sb_3__1_ sb_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_4__5__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_4__5__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_4__5__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_4__5__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_4__5__undriven_ccff_head),
		.chany_top_out(sb_4__5__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_4__5__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_4__5__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_4__5__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_4__5__undriven_ccff_tail));

	sb_3__1_ sb_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_4__6__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_4__6__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_4__6__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_4__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_4__6__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_4__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_4__6__undriven_ccff_head),
		.chany_top_out(sb_4__6__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_4__6__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_4__6__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_4__6__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_4__6__undriven_ccff_tail));

	sb_3__1_ sb_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_5__6__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_5__6__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_5__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_5__6__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_5__6__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_5__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_5__6__undriven_ccff_head),
		.chany_top_out(sb_5__6__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_5__6__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_5__6__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_5__6__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_5__6__undriven_ccff_tail));

	sb_5__0_ sb_5__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_5__0__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_36_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_36_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_37_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_37_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_38_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_38_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_39_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_39_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_40_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_40_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_41_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_41_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_42_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_42_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_43_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_43_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_44_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_44_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_45_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_45_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_46_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_46_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_47_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_47_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_48_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_48_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_49_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_49_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_50_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_50_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_51_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_51_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_52_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_52_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_53_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_53_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_54_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_54_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_55_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_55_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_56_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_56_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_57_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_57_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_58_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_58_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_59_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_59_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_60_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_60_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_61_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_61_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_62_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_62_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_63_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_63_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_64_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_64_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_65_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_65_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_66_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_66_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_67_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_67_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_68_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_68_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_69_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_69_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_70_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_70_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_out_71_(sb_5__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_out_71_),
		.chanx_right_in(sb_5__0__undriven_chanx_right_in[0:149]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_5__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(sb_5__0__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_5__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_5__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_5__0__undriven_ccff_head),
		.chany_top_out(sb_5__0__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_5__0__undriven_chanx_right_out[0:149]),
		.chanx_left_out(sb_5__0__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_5__0__undriven_ccff_tail));

	sb_5__1_ sb_5__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_5__1__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(sb_5__1__undriven_chany_bottom_in[0:149]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_36_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_36_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_37_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_37_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_38_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_38_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_39_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_39_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_40_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_40_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_41_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_41_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_42_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_42_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_43_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_43_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_44_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_44_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_45_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_45_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_46_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_46_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_47_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_47_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_48_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_48_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_49_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_49_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_50_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_50_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_51_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_51_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_52_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_52_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_53_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_53_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_54_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_54_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_55_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_55_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_56_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_56_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_57_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_57_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_58_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_58_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_59_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_59_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_60_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_60_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_61_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_61_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_62_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_62_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_63_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_63_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_64_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_64_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_65_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_65_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_66_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_66_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_67_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_67_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_68_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_68_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_69_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_69_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_70_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_70_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_71_(sb_5__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_out_71_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_5__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_5__1__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_5__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_5__1__undriven_ccff_head),
		.chany_top_out(sb_5__1__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_5__1__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_5__1__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_5__1__undriven_ccff_tail));

	sb_6__0_ sb_6__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_6__0__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_(sb_6__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_),
		.chanx_right_in(sb_6__0__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_6__0__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_6__0__undriven_right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(sb_6__0__undriven_chanx_left_in[0:149]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_6__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_6__0__undriven_ccff_head),
		.chany_top_out(sb_6__0__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_6__0__undriven_chanx_right_out[0:149]),
		.chanx_left_out(sb_6__0__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_6__0__undriven_ccff_tail));

	sb_6__1_ sb_6__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_6__1__undriven_chany_top_in[0:149]),
		.chanx_right_in(sb_6__1__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_6__1__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_6__1__undriven_chany_bottom_in[0:149]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_0_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_1_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_2_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_3_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_4_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_5_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_6_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_7_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_8_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_9_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_10_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_11_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_12_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_13_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_14_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_15_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_16_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_17_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_18_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_19_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_20_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_21_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_22_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_23_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_24_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_25_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_26_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_27_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_28_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_29_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_30_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_31_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_32_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_33_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_34_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_35_(sb_6__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_out_35_),
		.ccff_head(sb_6__1__undriven_ccff_head),
		.chany_top_out(sb_6__1__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_6__1__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_6__1__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_6__1__undriven_ccff_tail));

	sb_6__2_ sb_6__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_6__2__undriven_chany_top_in[0:149]),
		.chanx_right_in(sb_6__2__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_6__2__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_6__2__undriven_chany_bottom_in[0:149]),
		.ccff_head(sb_6__2__undriven_ccff_head),
		.chany_top_out(sb_6__2__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_6__2__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_6__2__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_6__2__undriven_ccff_tail));

	sb_6__2_ sb_6__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_6__3__undriven_chany_top_in[0:149]),
		.chanx_right_in(sb_6__3__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_6__3__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_6__3__undriven_chany_bottom_in[0:149]),
		.ccff_head(sb_6__3__undriven_ccff_head),
		.chany_top_out(sb_6__3__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_6__3__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_6__3__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_6__3__undriven_ccff_tail));

	sb_6__2_ sb_6__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_6__4__undriven_chany_top_in[0:149]),
		.chanx_right_in(sb_6__4__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_6__4__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_6__4__undriven_chany_bottom_in[0:149]),
		.ccff_head(sb_6__4__undriven_ccff_head),
		.chany_top_out(sb_6__4__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_6__4__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_6__4__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_6__4__undriven_ccff_tail));

	sb_6__2_ sb_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_6__5__undriven_chany_top_in[0:149]),
		.chanx_right_in(sb_6__5__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_6__5__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_6__5__undriven_chany_bottom_in[0:149]),
		.ccff_head(sb_6__5__undriven_ccff_head),
		.chany_top_out(sb_6__5__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_6__5__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_6__5__undriven_chany_bottom_out[0:149]),
		.ccff_tail(sb_6__5__undriven_ccff_tail));

	sb_6__6_ sb_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_6__6__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_6__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(sb_6__6__undriven_chanx_right_in[0:149]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_6__6__undriven_right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(sb_6__6__undriven_chany_bottom_in[0:149]),
		.chanx_left_in(sb_6__6__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_6__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_6__6__undriven_ccff_head),
		.chany_top_out(sb_6__6__undriven_chany_top_out[0:149]),
		.chanx_right_out(sb_6__6__undriven_chanx_right_out[0:149]),
		.chany_bottom_out(sb_6__6__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_6__6__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_6__6__undriven_ccff_tail));

	sb_7__0_ sb_7__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_7__0__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__0__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__0__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(sb_7__0__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_7__0__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__0__undriven_left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_7__0__undriven_ccff_head),
		.chany_top_out(sb_7__0__undriven_chany_top_out[0:149]),
		.chanx_left_out(sb_7__0__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_7__0__undriven_ccff_tail));

	sb_7__1_ sb_7__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_7__1__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__1__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__1__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_7__1__undriven_chany_bottom_in[0:149]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__1__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__1__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_7__1__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_7__1__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_7__1__undriven_ccff_head),
		.chany_top_out(sb_7__1__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_7__1__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_7__1__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_7__1__undriven_ccff_tail));

	sb_7__1_ sb_7__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_7__2__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__2__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__2__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_7__2__undriven_chany_bottom_in[0:149]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__2__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__2__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_7__2__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_7__2__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_7__2__undriven_ccff_head),
		.chany_top_out(sb_7__2__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_7__2__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_7__2__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_7__2__undriven_ccff_tail));

	sb_7__1_ sb_7__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_7__3__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__3__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__3__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_7__3__undriven_chany_bottom_in[0:149]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__3__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__3__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_7__3__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_7__3__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_7__3__undriven_ccff_head),
		.chany_top_out(sb_7__3__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_7__3__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_7__3__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_7__3__undriven_ccff_tail));

	sb_7__1_ sb_7__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_7__4__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__4__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__4__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_7__4__undriven_chany_bottom_in[0:149]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__4__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__4__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_7__4__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_7__4__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_7__4__undriven_ccff_head),
		.chany_top_out(sb_7__4__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_7__4__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_7__4__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_7__4__undriven_ccff_tail));

	sb_7__1_ sb_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_7__5__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__5__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__5__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_7__5__undriven_chany_bottom_in[0:149]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__5__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__5__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_7__5__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_7__5__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_7__5__undriven_ccff_head),
		.chany_top_out(sb_7__5__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_7__5__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_7__5__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_7__5__undriven_ccff_tail));

	sb_7__1_ sb_7__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(sb_7__6__undriven_chany_top_in[0:149]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__6__undriven_top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__6__undriven_top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(sb_7__6__undriven_chany_bottom_in[0:149]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__6__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__6__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_7__6__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(sb_7__6__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(sb_7__6__undriven_ccff_head),
		.chany_top_out(sb_7__6__undriven_chany_top_out[0:149]),
		.chany_bottom_out(sb_7__6__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_7__6__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_7__6__undriven_ccff_tail));

	sb_7__7_ sb_7__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_7__7__undriven_chany_bottom_in[0:149]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__7__undriven_bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_7__7__undriven_bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(sb_7__7__undriven_chanx_left_in[0:149]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(sb_7__7__undriven_left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_7__7__undriven_ccff_head),
		.chany_bottom_out(sb_7__7__undriven_chany_bottom_out[0:149]),
		.chanx_left_out(sb_7__7__undriven_chanx_left_out[0:149]),
		.ccff_tail(sb_7__7__undriven_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_1__0__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_1__0__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_1__0__undriven_ccff_head),
		.chanx_left_out(cbx_1__0__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_1__0__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_1__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__undriven_ccff_tail));

	cbx_1__0_ cbx_3__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_3__0__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_3__0__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_3__0__undriven_ccff_head),
		.chanx_left_out(cbx_3__0__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_3__0__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_3__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_3__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_3__0__undriven_ccff_tail));

	cbx_1__0_ cbx_4__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_4__0__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_4__0__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_4__0__undriven_ccff_head),
		.chanx_left_out(cbx_4__0__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_4__0__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_4__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_4__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_4__0__undriven_ccff_tail));

	cbx_1__0_ cbx_5__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_5__0__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_5__0__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_5__0__undriven_ccff_head),
		.chanx_left_out(cbx_5__0__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_5__0__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_5__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_5__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_5__0__undriven_ccff_tail));

	cbx_1__0_ cbx_7__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_7__0__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_7__0__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_7__0__undriven_ccff_head),
		.chanx_left_out(cbx_7__0__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_7__0__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_7__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_7__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_7__0__undriven_ccff_tail));

	cbx_1__1_ cbx_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_1__1__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_1__1__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_1__1__undriven_ccff_head),
		.chanx_left_out(cbx_1__1__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_1__1__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_1__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_1__1__undriven_ccff_tail));

	cbx_1__1_ cbx_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_1__2__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_1__2__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_1__2__undriven_ccff_head),
		.chanx_left_out(cbx_1__2__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_1__2__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_1__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_1__2__undriven_ccff_tail));

	cbx_1__1_ cbx_1__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_1__3__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_1__3__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_1__3__undriven_ccff_head),
		.chanx_left_out(cbx_1__3__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_1__3__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_1__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_1__3__undriven_ccff_tail));

	cbx_1__1_ cbx_1__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_1__4__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_1__4__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_1__4__undriven_ccff_head),
		.chanx_left_out(cbx_1__4__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_1__4__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_1__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_1__4__undriven_ccff_tail));

	cbx_1__1_ cbx_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_1__5__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_1__5__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_1__5__undriven_ccff_head),
		.chanx_left_out(cbx_1__5__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_1__5__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_1__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_1__5__undriven_ccff_tail));

	cbx_1__1_ cbx_1__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_1__6__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_1__6__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_1__6__undriven_ccff_head),
		.chanx_left_out(cbx_1__6__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_1__6__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_1__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_1__6__undriven_ccff_tail));

	cbx_1__1_ cbx_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_3__1__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_3__1__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_3__1__undriven_ccff_head),
		.chanx_left_out(cbx_3__1__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_3__1__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_3__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_3__1__undriven_ccff_tail));

	cbx_1__1_ cbx_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_3__2__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_3__2__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_3__2__undriven_ccff_head),
		.chanx_left_out(cbx_3__2__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_3__2__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_3__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_3__2__undriven_ccff_tail));

	cbx_1__1_ cbx_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_3__3__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_3__3__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_3__3__undriven_ccff_head),
		.chanx_left_out(cbx_3__3__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_3__3__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_3__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_3__3__undriven_ccff_tail));

	cbx_1__1_ cbx_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_3__4__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_3__4__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_3__4__undriven_ccff_head),
		.chanx_left_out(cbx_3__4__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_3__4__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_3__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_3__4__undriven_ccff_tail));

	cbx_1__1_ cbx_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_3__5__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_3__5__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_3__5__undriven_ccff_head),
		.chanx_left_out(cbx_3__5__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_3__5__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_3__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_3__5__undriven_ccff_tail));

	cbx_1__1_ cbx_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_3__6__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_3__6__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_3__6__undriven_ccff_head),
		.chanx_left_out(cbx_3__6__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_3__6__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_3__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_3__6__undriven_ccff_tail));

	cbx_1__1_ cbx_4__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_4__1__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_4__1__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_4__1__undriven_ccff_head),
		.chanx_left_out(cbx_4__1__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_4__1__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_4__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_4__1__undriven_ccff_tail));

	cbx_1__1_ cbx_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_4__2__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_4__2__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_4__2__undriven_ccff_head),
		.chanx_left_out(cbx_4__2__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_4__2__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_4__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_4__2__undriven_ccff_tail));

	cbx_1__1_ cbx_4__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_4__3__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_4__3__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_4__3__undriven_ccff_head),
		.chanx_left_out(cbx_4__3__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_4__3__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_4__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_4__3__undriven_ccff_tail));

	cbx_1__1_ cbx_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_4__4__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_4__4__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_4__4__undriven_ccff_head),
		.chanx_left_out(cbx_4__4__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_4__4__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_4__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_4__4__undriven_ccff_tail));

	cbx_1__1_ cbx_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_4__5__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_4__5__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_4__5__undriven_ccff_head),
		.chanx_left_out(cbx_4__5__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_4__5__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_4__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_4__5__undriven_ccff_tail));

	cbx_1__1_ cbx_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_4__6__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_4__6__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_4__6__undriven_ccff_head),
		.chanx_left_out(cbx_4__6__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_4__6__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_4__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_4__6__undriven_ccff_tail));

	cbx_1__1_ cbx_5__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_5__1__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_5__1__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_5__1__undriven_ccff_head),
		.chanx_left_out(cbx_5__1__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_5__1__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_5__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_5__1__undriven_ccff_tail));

	cbx_1__1_ cbx_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_5__2__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_5__2__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_5__2__undriven_ccff_head),
		.chanx_left_out(cbx_5__2__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_5__2__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_5__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_5__2__undriven_ccff_tail));

	cbx_1__1_ cbx_5__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_5__3__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_5__3__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_5__3__undriven_ccff_head),
		.chanx_left_out(cbx_5__3__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_5__3__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_5__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_5__3__undriven_ccff_tail));

	cbx_1__1_ cbx_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_5__4__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_5__4__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_5__4__undriven_ccff_head),
		.chanx_left_out(cbx_5__4__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_5__4__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_5__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_5__4__undriven_ccff_tail));

	cbx_1__1_ cbx_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_5__5__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_5__5__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_5__5__undriven_ccff_head),
		.chanx_left_out(cbx_5__5__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_5__5__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_5__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_5__5__undriven_ccff_tail));

	cbx_1__1_ cbx_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_5__6__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_5__6__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_5__6__undriven_ccff_head),
		.chanx_left_out(cbx_5__6__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_5__6__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_5__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_5__6__undriven_ccff_tail));

	cbx_1__1_ cbx_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_6__6__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_6__6__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_6__6__undriven_ccff_head),
		.chanx_left_out(cbx_6__6__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_6__6__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_6__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_6__6__undriven_ccff_tail));

	cbx_1__1_ cbx_7__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_7__1__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_7__1__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_7__1__undriven_ccff_head),
		.chanx_left_out(cbx_7__1__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_7__1__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_7__1__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_7__1__undriven_ccff_tail));

	cbx_1__1_ cbx_7__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_7__2__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_7__2__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_7__2__undriven_ccff_head),
		.chanx_left_out(cbx_7__2__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_7__2__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_7__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_7__2__undriven_ccff_tail));

	cbx_1__1_ cbx_7__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_7__3__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_7__3__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_7__3__undriven_ccff_head),
		.chanx_left_out(cbx_7__3__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_7__3__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_7__3__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_7__3__undriven_ccff_tail));

	cbx_1__1_ cbx_7__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_7__4__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_7__4__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_7__4__undriven_ccff_head),
		.chanx_left_out(cbx_7__4__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_7__4__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_7__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_7__4__undriven_ccff_tail));

	cbx_1__1_ cbx_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_7__5__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_7__5__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_7__5__undriven_ccff_head),
		.chanx_left_out(cbx_7__5__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_7__5__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_7__5__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_7__5__undriven_ccff_tail));

	cbx_1__1_ cbx_7__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_7__6__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_7__6__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_7__6__undriven_ccff_head),
		.chanx_left_out(cbx_7__6__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_7__6__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_7__6__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_7__6__undriven_ccff_tail));

	cbx_1__7_ cbx_1__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_1__7__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_1__7__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_1__7__undriven_ccff_head),
		.chanx_left_out(cbx_1__7__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_1__7__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__7__undriven_ccff_tail));

	cbx_1__7_ cbx_2__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_2__7__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_2__7__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_2__7__undriven_ccff_head),
		.chanx_left_out(cbx_2__7__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_2__7__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_2__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_2__7__undriven_ccff_tail));

	cbx_1__7_ cbx_3__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_3__7__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_3__7__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_3__7__undriven_ccff_head),
		.chanx_left_out(cbx_3__7__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_3__7__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_3__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_3__7__undriven_ccff_tail));

	cbx_1__7_ cbx_4__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_4__7__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_4__7__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_4__7__undriven_ccff_head),
		.chanx_left_out(cbx_4__7__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_4__7__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_4__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_4__7__undriven_ccff_tail));

	cbx_1__7_ cbx_5__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_5__7__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_5__7__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_5__7__undriven_ccff_head),
		.chanx_left_out(cbx_5__7__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_5__7__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_5__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_5__7__undriven_ccff_tail));

	cbx_1__7_ cbx_6__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_6__7__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_6__7__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_6__7__undriven_ccff_head),
		.chanx_left_out(cbx_6__7__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_6__7__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_6__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_6__7__undriven_ccff_tail));

	cbx_1__7_ cbx_7__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_7__7__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_7__7__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_7__7__undriven_ccff_head),
		.chanx_left_out(cbx_7__7__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_7__7__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_7__7__undriven_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_7__7__undriven_ccff_tail));

	cbx_2__0_ cbx_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_2__0__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_2__0__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_2__0__undriven_ccff_head),
		.chanx_left_out(cbx_2__0__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_2__0__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_(cbx_2__0__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_2__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_2__0__undriven_ccff_tail));

	cbx_2__2_ cbx_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_2__2__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_2__2__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_2__2__undriven_ccff_head),
		.chanx_left_out(cbx_2__2__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_2__2__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_(cbx_2__2__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_),
		.ccff_tail(cbx_2__2__undriven_ccff_tail));

	cbx_2__2_ cbx_2__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_2__4__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_2__4__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_2__4__undriven_ccff_head),
		.chanx_left_out(cbx_2__4__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_2__4__undriven_chanx_right_out[0:149]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_(cbx_2__4__undriven_top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_),
		.ccff_tail(cbx_2__4__undriven_ccff_tail));

	cbx_2__6_ cbx_2__6_ (
		.chanx_left_in(cbx_2__6__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_2__6__undriven_chanx_right_in[0:149]),
		.chanx_left_out(cbx_2__6__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_2__6__undriven_chanx_right_out[0:149]));

	cbx_6__0_ cbx_6__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_6__0__undriven_chanx_left_in[0:149]),
		.chanx_right_in(cbx_6__0__undriven_chanx_right_in[0:149]),
		.ccff_head(cbx_6__0__undriven_ccff_head),
		.chanx_left_out(cbx_6__0__undriven_chanx_left_out[0:149]),
		.chanx_right_out(cbx_6__0__undriven_chanx_right_out[0:149]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_6__0__undriven_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_6__0__undriven_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_0__1__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_0__1__undriven_chany_top_in[0:149]),
		.ccff_head(cby_0__1__undriven_ccff_head),
		.chany_bottom_out(cby_0__1__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_0__1__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__undriven_ccff_tail));

	cby_0__1_ cby_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_0__2__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_0__2__undriven_chany_top_in[0:149]),
		.ccff_head(cby_0__2__undriven_ccff_head),
		.chany_bottom_out(cby_0__2__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_0__2__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__2__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__2__undriven_ccff_tail));

	cby_0__1_ cby_0__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_0__3__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_0__3__undriven_chany_top_in[0:149]),
		.ccff_head(cby_0__3__undriven_ccff_head),
		.chany_bottom_out(cby_0__3__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_0__3__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__3__undriven_ccff_tail));

	cby_0__1_ cby_0__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_0__4__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_0__4__undriven_chany_top_in[0:149]),
		.ccff_head(cby_0__4__undriven_ccff_head),
		.chany_bottom_out(cby_0__4__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_0__4__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__4__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__4__undriven_ccff_tail));

	cby_0__1_ cby_0__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_0__5__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_0__5__undriven_chany_top_in[0:149]),
		.ccff_head(cby_0__5__undriven_ccff_head),
		.chany_bottom_out(cby_0__5__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_0__5__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__5__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__5__undriven_ccff_tail));

	cby_0__1_ cby_0__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_0__6__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_0__6__undriven_chany_top_in[0:149]),
		.ccff_head(cby_0__6__undriven_ccff_head),
		.chany_bottom_out(cby_0__6__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_0__6__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__6__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__6__undriven_ccff_tail));

	cby_0__1_ cby_0__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_0__7__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_0__7__undriven_chany_top_in[0:149]),
		.ccff_head(cby_0__7__undriven_ccff_head),
		.chany_bottom_out(cby_0__7__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_0__7__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__7__undriven_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__7__undriven_ccff_tail));

	cby_1__1_ cby_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_1__1__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_1__1__undriven_chany_top_in[0:149]),
		.ccff_head(cby_1__1__undriven_ccff_head),
		.chany_bottom_out(cby_1__1__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_1__1__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_1__1__undriven_ccff_tail));

	cby_1__1_ cby_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_1__2__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_1__2__undriven_chany_top_in[0:149]),
		.ccff_head(cby_1__2__undriven_ccff_head),
		.chany_bottom_out(cby_1__2__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_1__2__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_1__2__undriven_ccff_tail));

	cby_1__1_ cby_1__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_1__3__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_1__3__undriven_chany_top_in[0:149]),
		.ccff_head(cby_1__3__undriven_ccff_head),
		.chany_bottom_out(cby_1__3__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_1__3__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_1__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_1__3__undriven_ccff_tail));

	cby_1__1_ cby_1__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_1__4__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_1__4__undriven_chany_top_in[0:149]),
		.ccff_head(cby_1__4__undriven_ccff_head),
		.chany_bottom_out(cby_1__4__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_1__4__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_1__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_1__4__undriven_ccff_tail));

	cby_1__1_ cby_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_1__5__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_1__5__undriven_chany_top_in[0:149]),
		.ccff_head(cby_1__5__undriven_ccff_head),
		.chany_bottom_out(cby_1__5__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_1__5__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_1__5__undriven_ccff_tail));

	cby_1__1_ cby_1__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_1__6__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_1__6__undriven_chany_top_in[0:149]),
		.ccff_head(cby_1__6__undriven_ccff_head),
		.chany_bottom_out(cby_1__6__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_1__6__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_1__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_1__6__undriven_ccff_tail));

	cby_1__1_ cby_1__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_1__7__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_1__7__undriven_chany_top_in[0:149]),
		.ccff_head(cby_1__7__undriven_ccff_head),
		.chany_bottom_out(cby_1__7__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_1__7__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_1__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_1__7__undriven_ccff_tail));

	cby_1__1_ cby_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_3__1__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_3__1__undriven_chany_top_in[0:149]),
		.ccff_head(cby_3__1__undriven_ccff_head),
		.chany_bottom_out(cby_3__1__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_3__1__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_3__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_3__1__undriven_ccff_tail));

	cby_1__1_ cby_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_3__2__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_3__2__undriven_chany_top_in[0:149]),
		.ccff_head(cby_3__2__undriven_ccff_head),
		.chany_bottom_out(cby_3__2__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_3__2__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_3__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_3__2__undriven_ccff_tail));

	cby_1__1_ cby_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_3__3__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_3__3__undriven_chany_top_in[0:149]),
		.ccff_head(cby_3__3__undriven_ccff_head),
		.chany_bottom_out(cby_3__3__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_3__3__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_3__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_3__3__undriven_ccff_tail));

	cby_1__1_ cby_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_3__4__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_3__4__undriven_chany_top_in[0:149]),
		.ccff_head(cby_3__4__undriven_ccff_head),
		.chany_bottom_out(cby_3__4__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_3__4__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_3__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_3__4__undriven_ccff_tail));

	cby_1__1_ cby_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_3__5__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_3__5__undriven_chany_top_in[0:149]),
		.ccff_head(cby_3__5__undriven_ccff_head),
		.chany_bottom_out(cby_3__5__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_3__5__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_3__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_3__5__undriven_ccff_tail));

	cby_1__1_ cby_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_3__6__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_3__6__undriven_chany_top_in[0:149]),
		.ccff_head(cby_3__6__undriven_ccff_head),
		.chany_bottom_out(cby_3__6__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_3__6__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_3__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_3__6__undriven_ccff_tail));

	cby_1__1_ cby_3__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_3__7__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_3__7__undriven_chany_top_in[0:149]),
		.ccff_head(cby_3__7__undriven_ccff_head),
		.chany_bottom_out(cby_3__7__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_3__7__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_3__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_3__7__undriven_ccff_tail));

	cby_1__1_ cby_4__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_4__1__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_4__1__undriven_chany_top_in[0:149]),
		.ccff_head(cby_4__1__undriven_ccff_head),
		.chany_bottom_out(cby_4__1__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_4__1__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_4__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_4__1__undriven_ccff_tail));

	cby_1__1_ cby_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_4__2__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_4__2__undriven_chany_top_in[0:149]),
		.ccff_head(cby_4__2__undriven_ccff_head),
		.chany_bottom_out(cby_4__2__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_4__2__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_4__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_4__2__undriven_ccff_tail));

	cby_1__1_ cby_4__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_4__3__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_4__3__undriven_chany_top_in[0:149]),
		.ccff_head(cby_4__3__undriven_ccff_head),
		.chany_bottom_out(cby_4__3__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_4__3__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_4__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_4__3__undriven_ccff_tail));

	cby_1__1_ cby_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_4__4__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_4__4__undriven_chany_top_in[0:149]),
		.ccff_head(cby_4__4__undriven_ccff_head),
		.chany_bottom_out(cby_4__4__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_4__4__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_4__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_4__4__undriven_ccff_tail));

	cby_1__1_ cby_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_4__5__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_4__5__undriven_chany_top_in[0:149]),
		.ccff_head(cby_4__5__undriven_ccff_head),
		.chany_bottom_out(cby_4__5__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_4__5__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_4__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_4__5__undriven_ccff_tail));

	cby_1__1_ cby_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_4__6__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_4__6__undriven_chany_top_in[0:149]),
		.ccff_head(cby_4__6__undriven_ccff_head),
		.chany_bottom_out(cby_4__6__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_4__6__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_4__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_4__6__undriven_ccff_tail));

	cby_1__1_ cby_4__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_4__7__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_4__7__undriven_chany_top_in[0:149]),
		.ccff_head(cby_4__7__undriven_ccff_head),
		.chany_bottom_out(cby_4__7__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_4__7__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_4__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_4__7__undriven_ccff_tail));

	cby_1__1_ cby_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_5__2__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_5__2__undriven_chany_top_in[0:149]),
		.ccff_head(cby_5__2__undriven_ccff_head),
		.chany_bottom_out(cby_5__2__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_5__2__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_5__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_5__2__undriven_ccff_tail));

	cby_1__1_ cby_5__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_5__3__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_5__3__undriven_chany_top_in[0:149]),
		.ccff_head(cby_5__3__undriven_ccff_head),
		.chany_bottom_out(cby_5__3__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_5__3__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_5__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_5__3__undriven_ccff_tail));

	cby_1__1_ cby_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_5__4__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_5__4__undriven_chany_top_in[0:149]),
		.ccff_head(cby_5__4__undriven_ccff_head),
		.chany_bottom_out(cby_5__4__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_5__4__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_5__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_5__4__undriven_ccff_tail));

	cby_1__1_ cby_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_5__5__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_5__5__undriven_chany_top_in[0:149]),
		.ccff_head(cby_5__5__undriven_ccff_head),
		.chany_bottom_out(cby_5__5__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_5__5__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_5__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_5__5__undriven_ccff_tail));

	cby_1__1_ cby_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_5__6__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_5__6__undriven_chany_top_in[0:149]),
		.ccff_head(cby_5__6__undriven_ccff_head),
		.chany_bottom_out(cby_5__6__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_5__6__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_5__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_5__6__undriven_ccff_tail));

	cby_1__1_ cby_5__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_5__7__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_5__7__undriven_chany_top_in[0:149]),
		.ccff_head(cby_5__7__undriven_ccff_head),
		.chany_bottom_out(cby_5__7__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_5__7__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_5__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_5__7__undriven_ccff_tail));

	cby_1__1_ cby_6__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_6__7__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_6__7__undriven_chany_top_in[0:149]),
		.ccff_head(cby_6__7__undriven_ccff_head),
		.chany_bottom_out(cby_6__7__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_6__7__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_6__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_6__7__undriven_ccff_tail));

	cby_2__1_ cby_2__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_2__1__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_2__1__undriven_chany_top_in[0:149]),
		.ccff_head(cby_2__1__undriven_ccff_head),
		.chany_bottom_out(cby_2__1__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_2__1__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_2__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_2__1__undriven_ccff_tail));

	cby_2__1_ cby_2__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_2__3__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_2__3__undriven_chany_top_in[0:149]),
		.ccff_head(cby_2__3__undriven_ccff_head),
		.chany_bottom_out(cby_2__3__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_2__3__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_2__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_2__3__undriven_ccff_tail));

	cby_2__1_ cby_2__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_2__5__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_2__5__undriven_chany_top_in[0:149]),
		.ccff_head(cby_2__5__undriven_ccff_head),
		.chany_bottom_out(cby_2__5__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_2__5__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_2__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_2__5__undriven_ccff_tail));

	cby_2__2_ cby_2__2_ (
		.chany_bottom_in(cby_2__2__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_2__2__undriven_chany_top_in[0:149]),
		.chany_bottom_out(cby_2__2__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_2__2__undriven_chany_top_out[0:149]));

	cby_2__2_ cby_2__4_ (
		.chany_bottom_in(cby_2__4__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_2__4__undriven_chany_top_in[0:149]),
		.chany_bottom_out(cby_2__4__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_2__4__undriven_chany_top_out[0:149]));

	cby_2__2_ cby_2__6_ (
		.chany_bottom_in(cby_2__6__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_2__6__undriven_chany_top_in[0:149]),
		.chany_bottom_out(cby_2__6__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_2__6__undriven_chany_top_out[0:149]));

	cby_2__2_ cby_2__7_ (
		.chany_bottom_in(cby_2__7__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_2__7__undriven_chany_top_in[0:149]),
		.chany_bottom_out(cby_2__7__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_2__7__undriven_chany_top_out[0:149]));

	cby_2__2_ cby_6__2_ (
		.chany_bottom_in(cby_6__2__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_6__2__undriven_chany_top_in[0:149]),
		.chany_bottom_out(cby_6__2__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_6__2__undriven_chany_top_out[0:149]));

	cby_2__2_ cby_6__3_ (
		.chany_bottom_in(cby_6__3__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_6__3__undriven_chany_top_in[0:149]),
		.chany_bottom_out(cby_6__3__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_6__3__undriven_chany_top_out[0:149]));

	cby_2__2_ cby_6__4_ (
		.chany_bottom_in(cby_6__4__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_6__4__undriven_chany_top_in[0:149]),
		.chany_bottom_out(cby_6__4__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_6__4__undriven_chany_top_out[0:149]));

	cby_2__2_ cby_6__5_ (
		.chany_bottom_in(cby_6__5__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_6__5__undriven_chany_top_in[0:149]),
		.chany_bottom_out(cby_6__5__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_6__5__undriven_chany_top_out[0:149]));

	cby_2__2_ cby_6__6_ (
		.chany_bottom_in(cby_6__6__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_6__6__undriven_chany_top_in[0:149]),
		.chany_bottom_out(cby_6__6__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_6__6__undriven_chany_top_out[0:149]));

	cby_5__1_ cby_5__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_5__1__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_5__1__undriven_chany_top_in[0:149]),
		.ccff_head(cby_5__1__undriven_ccff_head),
		.chany_bottom_out(cby_5__1__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_5__1__undriven_chany_top_out[0:149]),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_0_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_1_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_2_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_3_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_4_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_5_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_6_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_7_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_8_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_9_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_10_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_11_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_12_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_13_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_14_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_15_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_16_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_17_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_18_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_19_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_20_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_21_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_22_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_23_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_24_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_25_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_26_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_27_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_28_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_29_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_30_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_31_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_32_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_33_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_34_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_b_35_(cby_5__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_b_35_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_5__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_5__1__undriven_ccff_tail));

	cby_6__1_ cby_6__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_6__1__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_6__1__undriven_chany_top_in[0:149]),
		.ccff_head(cby_6__1__undriven_ccff_head),
		.chany_bottom_out(cby_6__1__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_6__1__undriven_chany_top_out[0:149]),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_0_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_1_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_2_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_3_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_4_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_5_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_6_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_7_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_8_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_9_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_10_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_11_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_12_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_13_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_14_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_15_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_16_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_17_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_18_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_19_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_20_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_21_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_22_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_23_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_24_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_25_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_26_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_27_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_28_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_29_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_30_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_31_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_32_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_33_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_34_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_35_(cby_6__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_a_35_),
		.ccff_tail(cby_6__1__undriven_ccff_tail));

	cby_7__1_ cby_7__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_7__1__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_7__1__undriven_chany_top_in[0:149]),
		.ccff_head(cby_7__1__undriven_ccff_head),
		.chany_bottom_out(cby_7__1__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_7__1__undriven_chany_top_out[0:149]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_7__1__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_7__1__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_7__1__undriven_ccff_tail));

	cby_7__1_ cby_7__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_7__2__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_7__2__undriven_chany_top_in[0:149]),
		.ccff_head(cby_7__2__undriven_ccff_head),
		.chany_bottom_out(cby_7__2__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_7__2__undriven_chany_top_out[0:149]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_7__2__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_7__2__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_7__2__undriven_ccff_tail));

	cby_7__1_ cby_7__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_7__3__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_7__3__undriven_chany_top_in[0:149]),
		.ccff_head(cby_7__3__undriven_ccff_head),
		.chany_bottom_out(cby_7__3__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_7__3__undriven_chany_top_out[0:149]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_7__3__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_7__3__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_7__3__undriven_ccff_tail));

	cby_7__1_ cby_7__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_7__4__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_7__4__undriven_chany_top_in[0:149]),
		.ccff_head(cby_7__4__undriven_ccff_head),
		.chany_bottom_out(cby_7__4__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_7__4__undriven_chany_top_out[0:149]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_7__4__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_7__4__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_7__4__undriven_ccff_tail));

	cby_7__1_ cby_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_7__5__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_7__5__undriven_chany_top_in[0:149]),
		.ccff_head(cby_7__5__undriven_ccff_head),
		.chany_bottom_out(cby_7__5__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_7__5__undriven_chany_top_out[0:149]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_7__5__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_7__5__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_7__5__undriven_ccff_tail));

	cby_7__1_ cby_7__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_7__6__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_7__6__undriven_chany_top_in[0:149]),
		.ccff_head(cby_7__6__undriven_ccff_head),
		.chany_bottom_out(cby_7__6__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_7__6__undriven_chany_top_out[0:149]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_7__6__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_7__6__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_7__6__undriven_ccff_tail));

	cby_7__1_ cby_7__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_7__7__undriven_chany_bottom_in[0:149]),
		.chany_top_in(cby_7__7__undriven_chany_top_in[0:149]),
		.ccff_head(cby_7__7__undriven_ccff_head),
		.chany_bottom_out(cby_7__7__undriven_chany_bottom_out[0:149]),
		.chany_top_out(cby_7__7__undriven_chany_top_out[0:149]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_7__7__undriven_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_7__7__undriven_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_7__7__undriven_ccff_tail));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
`default_nettype wire




