//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[6][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Mon Jul  7 22:56:01 2025
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_6__0_ -----
module sb_6__0_(pReset,
                prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                chanx_left_in,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:149] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_;
//----- INPUT PORTS -----
input [0:149] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:149] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:149] chany_top_out;
//----- OUTPUT PORTS -----
output [0:149] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:149] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:7] mux_2level_tapbuf_size10_0_sram;
wire [0:7] mux_2level_tapbuf_size10_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_10_sram;
wire [0:7] mux_2level_tapbuf_size10_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_11_sram;
wire [0:7] mux_2level_tapbuf_size10_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_12_sram;
wire [0:7] mux_2level_tapbuf_size10_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_1_sram;
wire [0:7] mux_2level_tapbuf_size10_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_2_sram;
wire [0:7] mux_2level_tapbuf_size10_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_3_sram;
wire [0:7] mux_2level_tapbuf_size10_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_4_sram;
wire [0:7] mux_2level_tapbuf_size10_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_5_sram;
wire [0:7] mux_2level_tapbuf_size10_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_6_sram;
wire [0:7] mux_2level_tapbuf_size10_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_7_sram;
wire [0:7] mux_2level_tapbuf_size10_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_8_sram;
wire [0:7] mux_2level_tapbuf_size10_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_9_sram;
wire [0:7] mux_2level_tapbuf_size10_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size10_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size4_0_sram;
wire [0:5] mux_2level_tapbuf_size4_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_1_sram;
wire [0:5] mux_2level_tapbuf_size4_1_sram_inv;
wire [0:0] mux_2level_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_1_ccff_tail;
wire [0:5] mux_2level_tapbuf_size5_0_sram;
wire [0:5] mux_2level_tapbuf_size5_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_10_sram;
wire [0:5] mux_2level_tapbuf_size5_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_11_sram;
wire [0:5] mux_2level_tapbuf_size5_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_12_sram;
wire [0:5] mux_2level_tapbuf_size5_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_13_sram;
wire [0:5] mux_2level_tapbuf_size5_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_14_sram;
wire [0:5] mux_2level_tapbuf_size5_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_15_sram;
wire [0:5] mux_2level_tapbuf_size5_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_16_sram;
wire [0:5] mux_2level_tapbuf_size5_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_17_sram;
wire [0:5] mux_2level_tapbuf_size5_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_18_sram;
wire [0:5] mux_2level_tapbuf_size5_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_19_sram;
wire [0:5] mux_2level_tapbuf_size5_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_1_sram;
wire [0:5] mux_2level_tapbuf_size5_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_20_sram;
wire [0:5] mux_2level_tapbuf_size5_20_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_21_sram;
wire [0:5] mux_2level_tapbuf_size5_21_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_22_sram;
wire [0:5] mux_2level_tapbuf_size5_22_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_23_sram;
wire [0:5] mux_2level_tapbuf_size5_23_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_24_sram;
wire [0:5] mux_2level_tapbuf_size5_24_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_25_sram;
wire [0:5] mux_2level_tapbuf_size5_25_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_26_sram;
wire [0:5] mux_2level_tapbuf_size5_26_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_27_sram;
wire [0:5] mux_2level_tapbuf_size5_27_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_28_sram;
wire [0:5] mux_2level_tapbuf_size5_28_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_29_sram;
wire [0:5] mux_2level_tapbuf_size5_29_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_2_sram;
wire [0:5] mux_2level_tapbuf_size5_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_30_sram;
wire [0:5] mux_2level_tapbuf_size5_30_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_31_sram;
wire [0:5] mux_2level_tapbuf_size5_31_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_32_sram;
wire [0:5] mux_2level_tapbuf_size5_32_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_33_sram;
wire [0:5] mux_2level_tapbuf_size5_33_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_34_sram;
wire [0:5] mux_2level_tapbuf_size5_34_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_35_sram;
wire [0:5] mux_2level_tapbuf_size5_35_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_36_sram;
wire [0:5] mux_2level_tapbuf_size5_36_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_37_sram;
wire [0:5] mux_2level_tapbuf_size5_37_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_38_sram;
wire [0:5] mux_2level_tapbuf_size5_38_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_39_sram;
wire [0:5] mux_2level_tapbuf_size5_39_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_3_sram;
wire [0:5] mux_2level_tapbuf_size5_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_40_sram;
wire [0:5] mux_2level_tapbuf_size5_40_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_41_sram;
wire [0:5] mux_2level_tapbuf_size5_41_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_42_sram;
wire [0:5] mux_2level_tapbuf_size5_42_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_43_sram;
wire [0:5] mux_2level_tapbuf_size5_43_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_44_sram;
wire [0:5] mux_2level_tapbuf_size5_44_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_45_sram;
wire [0:5] mux_2level_tapbuf_size5_45_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_46_sram;
wire [0:5] mux_2level_tapbuf_size5_46_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_47_sram;
wire [0:5] mux_2level_tapbuf_size5_47_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_48_sram;
wire [0:5] mux_2level_tapbuf_size5_48_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_49_sram;
wire [0:5] mux_2level_tapbuf_size5_49_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_4_sram;
wire [0:5] mux_2level_tapbuf_size5_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_50_sram;
wire [0:5] mux_2level_tapbuf_size5_50_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_51_sram;
wire [0:5] mux_2level_tapbuf_size5_51_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_52_sram;
wire [0:5] mux_2level_tapbuf_size5_52_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_53_sram;
wire [0:5] mux_2level_tapbuf_size5_53_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_54_sram;
wire [0:5] mux_2level_tapbuf_size5_54_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_55_sram;
wire [0:5] mux_2level_tapbuf_size5_55_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_56_sram;
wire [0:5] mux_2level_tapbuf_size5_56_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_57_sram;
wire [0:5] mux_2level_tapbuf_size5_57_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_58_sram;
wire [0:5] mux_2level_tapbuf_size5_58_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_5_sram;
wire [0:5] mux_2level_tapbuf_size5_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_6_sram;
wire [0:5] mux_2level_tapbuf_size5_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_7_sram;
wire [0:5] mux_2level_tapbuf_size5_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_8_sram;
wire [0:5] mux_2level_tapbuf_size5_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_9_sram;
wire [0:5] mux_2level_tapbuf_size5_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size6_0_sram;
wire [0:5] mux_2level_tapbuf_size6_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_10_sram;
wire [0:5] mux_2level_tapbuf_size6_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_11_sram;
wire [0:5] mux_2level_tapbuf_size6_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_12_sram;
wire [0:5] mux_2level_tapbuf_size6_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_13_sram;
wire [0:5] mux_2level_tapbuf_size6_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_14_sram;
wire [0:5] mux_2level_tapbuf_size6_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_15_sram;
wire [0:5] mux_2level_tapbuf_size6_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_16_sram;
wire [0:5] mux_2level_tapbuf_size6_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_17_sram;
wire [0:5] mux_2level_tapbuf_size6_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_18_sram;
wire [0:5] mux_2level_tapbuf_size6_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_19_sram;
wire [0:5] mux_2level_tapbuf_size6_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_1_sram;
wire [0:5] mux_2level_tapbuf_size6_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_20_sram;
wire [0:5] mux_2level_tapbuf_size6_20_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_21_sram;
wire [0:5] mux_2level_tapbuf_size6_21_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_22_sram;
wire [0:5] mux_2level_tapbuf_size6_22_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_23_sram;
wire [0:5] mux_2level_tapbuf_size6_23_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_24_sram;
wire [0:5] mux_2level_tapbuf_size6_24_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_25_sram;
wire [0:5] mux_2level_tapbuf_size6_25_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_26_sram;
wire [0:5] mux_2level_tapbuf_size6_26_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_27_sram;
wire [0:5] mux_2level_tapbuf_size6_27_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_28_sram;
wire [0:5] mux_2level_tapbuf_size6_28_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_29_sram;
wire [0:5] mux_2level_tapbuf_size6_29_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_2_sram;
wire [0:5] mux_2level_tapbuf_size6_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_30_sram;
wire [0:5] mux_2level_tapbuf_size6_30_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_31_sram;
wire [0:5] mux_2level_tapbuf_size6_31_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_32_sram;
wire [0:5] mux_2level_tapbuf_size6_32_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_33_sram;
wire [0:5] mux_2level_tapbuf_size6_33_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_34_sram;
wire [0:5] mux_2level_tapbuf_size6_34_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_35_sram;
wire [0:5] mux_2level_tapbuf_size6_35_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_36_sram;
wire [0:5] mux_2level_tapbuf_size6_36_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_37_sram;
wire [0:5] mux_2level_tapbuf_size6_37_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_38_sram;
wire [0:5] mux_2level_tapbuf_size6_38_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_39_sram;
wire [0:5] mux_2level_tapbuf_size6_39_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_3_sram;
wire [0:5] mux_2level_tapbuf_size6_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_40_sram;
wire [0:5] mux_2level_tapbuf_size6_40_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_41_sram;
wire [0:5] mux_2level_tapbuf_size6_41_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_42_sram;
wire [0:5] mux_2level_tapbuf_size6_42_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_43_sram;
wire [0:5] mux_2level_tapbuf_size6_43_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_44_sram;
wire [0:5] mux_2level_tapbuf_size6_44_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_45_sram;
wire [0:5] mux_2level_tapbuf_size6_45_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_46_sram;
wire [0:5] mux_2level_tapbuf_size6_46_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_47_sram;
wire [0:5] mux_2level_tapbuf_size6_47_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_48_sram;
wire [0:5] mux_2level_tapbuf_size6_48_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_49_sram;
wire [0:5] mux_2level_tapbuf_size6_49_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_4_sram;
wire [0:5] mux_2level_tapbuf_size6_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_50_sram;
wire [0:5] mux_2level_tapbuf_size6_50_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_51_sram;
wire [0:5] mux_2level_tapbuf_size6_51_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_52_sram;
wire [0:5] mux_2level_tapbuf_size6_52_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_53_sram;
wire [0:5] mux_2level_tapbuf_size6_53_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_54_sram;
wire [0:5] mux_2level_tapbuf_size6_54_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_55_sram;
wire [0:5] mux_2level_tapbuf_size6_55_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_56_sram;
wire [0:5] mux_2level_tapbuf_size6_56_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_57_sram;
wire [0:5] mux_2level_tapbuf_size6_57_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_58_sram;
wire [0:5] mux_2level_tapbuf_size6_58_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_59_sram;
wire [0:5] mux_2level_tapbuf_size6_59_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_5_sram;
wire [0:5] mux_2level_tapbuf_size6_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_60_sram;
wire [0:5] mux_2level_tapbuf_size6_60_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_61_sram;
wire [0:5] mux_2level_tapbuf_size6_61_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_62_sram;
wire [0:5] mux_2level_tapbuf_size6_62_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_63_sram;
wire [0:5] mux_2level_tapbuf_size6_63_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_64_sram;
wire [0:5] mux_2level_tapbuf_size6_64_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_65_sram;
wire [0:5] mux_2level_tapbuf_size6_65_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_66_sram;
wire [0:5] mux_2level_tapbuf_size6_66_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_67_sram;
wire [0:5] mux_2level_tapbuf_size6_67_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_68_sram;
wire [0:5] mux_2level_tapbuf_size6_68_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_69_sram;
wire [0:5] mux_2level_tapbuf_size6_69_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_6_sram;
wire [0:5] mux_2level_tapbuf_size6_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_70_sram;
wire [0:5] mux_2level_tapbuf_size6_70_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_71_sram;
wire [0:5] mux_2level_tapbuf_size6_71_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_72_sram;
wire [0:5] mux_2level_tapbuf_size6_72_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_73_sram;
wire [0:5] mux_2level_tapbuf_size6_73_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_74_sram;
wire [0:5] mux_2level_tapbuf_size6_74_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_75_sram;
wire [0:5] mux_2level_tapbuf_size6_75_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_76_sram;
wire [0:5] mux_2level_tapbuf_size6_76_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_77_sram;
wire [0:5] mux_2level_tapbuf_size6_77_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_78_sram;
wire [0:5] mux_2level_tapbuf_size6_78_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_79_sram;
wire [0:5] mux_2level_tapbuf_size6_79_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_7_sram;
wire [0:5] mux_2level_tapbuf_size6_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_80_sram;
wire [0:5] mux_2level_tapbuf_size6_80_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_81_sram;
wire [0:5] mux_2level_tapbuf_size6_81_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_82_sram;
wire [0:5] mux_2level_tapbuf_size6_82_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_83_sram;
wire [0:5] mux_2level_tapbuf_size6_83_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_84_sram;
wire [0:5] mux_2level_tapbuf_size6_84_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_85_sram;
wire [0:5] mux_2level_tapbuf_size6_85_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_86_sram;
wire [0:5] mux_2level_tapbuf_size6_86_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_8_sram;
wire [0:5] mux_2level_tapbuf_size6_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_9_sram;
wire [0:5] mux_2level_tapbuf_size6_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_79_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_80_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_81_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_82_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_83_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_84_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_85_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_86_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size7_0_sram;
wire [0:5] mux_2level_tapbuf_size7_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_1_sram;
wire [0:5] mux_2level_tapbuf_size7_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_2_sram;
wire [0:5] mux_2level_tapbuf_size7_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_3_sram;
wire [0:5] mux_2level_tapbuf_size7_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_4_sram;
wire [0:5] mux_2level_tapbuf_size7_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_5_sram;
wire [0:5] mux_2level_tapbuf_size7_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_6_sram;
wire [0:5] mux_2level_tapbuf_size7_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_7_sram;
wire [0:5] mux_2level_tapbuf_size7_7_sram_inv;
wire [0:0] mux_2level_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_6_ccff_tail;
wire [0:5] mux_2level_tapbuf_size8_0_sram;
wire [0:5] mux_2level_tapbuf_size8_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_10_sram;
wire [0:5] mux_2level_tapbuf_size8_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_11_sram;
wire [0:5] mux_2level_tapbuf_size8_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_12_sram;
wire [0:5] mux_2level_tapbuf_size8_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_13_sram;
wire [0:5] mux_2level_tapbuf_size8_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_14_sram;
wire [0:5] mux_2level_tapbuf_size8_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_15_sram;
wire [0:5] mux_2level_tapbuf_size8_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_16_sram;
wire [0:5] mux_2level_tapbuf_size8_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_17_sram;
wire [0:5] mux_2level_tapbuf_size8_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_18_sram;
wire [0:5] mux_2level_tapbuf_size8_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_19_sram;
wire [0:5] mux_2level_tapbuf_size8_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_1_sram;
wire [0:5] mux_2level_tapbuf_size8_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_20_sram;
wire [0:5] mux_2level_tapbuf_size8_20_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_21_sram;
wire [0:5] mux_2level_tapbuf_size8_21_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_22_sram;
wire [0:5] mux_2level_tapbuf_size8_22_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_23_sram;
wire [0:5] mux_2level_tapbuf_size8_23_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_24_sram;
wire [0:5] mux_2level_tapbuf_size8_24_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_25_sram;
wire [0:5] mux_2level_tapbuf_size8_25_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_26_sram;
wire [0:5] mux_2level_tapbuf_size8_26_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_27_sram;
wire [0:5] mux_2level_tapbuf_size8_27_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_28_sram;
wire [0:5] mux_2level_tapbuf_size8_28_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_29_sram;
wire [0:5] mux_2level_tapbuf_size8_29_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_2_sram;
wire [0:5] mux_2level_tapbuf_size8_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_3_sram;
wire [0:5] mux_2level_tapbuf_size8_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_4_sram;
wire [0:5] mux_2level_tapbuf_size8_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_5_sram;
wire [0:5] mux_2level_tapbuf_size8_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_6_sram;
wire [0:5] mux_2level_tapbuf_size8_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_7_sram;
wire [0:5] mux_2level_tapbuf_size8_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_8_sram;
wire [0:5] mux_2level_tapbuf_size8_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_9_sram;
wire [0:5] mux_2level_tapbuf_size8_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size8_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_9_ccff_tail;
wire [0:7] mux_2level_tapbuf_size9_0_sram;
wire [0:7] mux_2level_tapbuf_size9_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_10_sram;
wire [0:7] mux_2level_tapbuf_size9_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_11_sram;
wire [0:7] mux_2level_tapbuf_size9_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_12_sram;
wire [0:7] mux_2level_tapbuf_size9_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_13_sram;
wire [0:7] mux_2level_tapbuf_size9_13_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_14_sram;
wire [0:7] mux_2level_tapbuf_size9_14_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_15_sram;
wire [0:7] mux_2level_tapbuf_size9_15_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_16_sram;
wire [0:7] mux_2level_tapbuf_size9_16_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_17_sram;
wire [0:7] mux_2level_tapbuf_size9_17_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_18_sram;
wire [0:7] mux_2level_tapbuf_size9_18_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_19_sram;
wire [0:7] mux_2level_tapbuf_size9_19_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_1_sram;
wire [0:7] mux_2level_tapbuf_size9_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_20_sram;
wire [0:7] mux_2level_tapbuf_size9_20_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_21_sram;
wire [0:7] mux_2level_tapbuf_size9_21_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_22_sram;
wire [0:7] mux_2level_tapbuf_size9_22_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_23_sram;
wire [0:7] mux_2level_tapbuf_size9_23_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_24_sram;
wire [0:7] mux_2level_tapbuf_size9_24_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_25_sram;
wire [0:7] mux_2level_tapbuf_size9_25_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_26_sram;
wire [0:7] mux_2level_tapbuf_size9_26_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_2_sram;
wire [0:7] mux_2level_tapbuf_size9_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_3_sram;
wire [0:7] mux_2level_tapbuf_size9_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_4_sram;
wire [0:7] mux_2level_tapbuf_size9_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_5_sram;
wire [0:7] mux_2level_tapbuf_size9_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_6_sram;
wire [0:7] mux_2level_tapbuf_size9_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_7_sram;
wire [0:7] mux_2level_tapbuf_size9_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_8_sram;
wire [0:7] mux_2level_tapbuf_size9_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_9_sram;
wire [0:7] mux_2level_tapbuf_size9_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size9_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[2] = chanx_right_in[1];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[6] = chanx_right_in[5];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[10] = chanx_right_in[9];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[83] = chanx_right_in[82];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[87] = chanx_right_in[86];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[91] = chanx_right_in[90];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[95] = chanx_right_in[94];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[97] = chanx_right_in[96];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[98] = chanx_right_in[97];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[99] = chanx_right_in[98];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[101] = chanx_right_in[100];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[102] = chanx_right_in[101];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[103] = chanx_right_in[102];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[105] = chanx_right_in[104];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[106] = chanx_right_in[105];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[107] = chanx_right_in[106];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[109] = chanx_right_in[108];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[110] = chanx_right_in[109];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[111] = chanx_right_in[110];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[113] = chanx_right_in[112];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[114] = chanx_right_in[113];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[115] = chanx_right_in[114];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[117] = chanx_right_in[116];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[118] = chanx_right_in[117];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[119] = chanx_right_in[118];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[121] = chanx_right_in[120];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[122] = chanx_right_in[121];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[123] = chanx_right_in[122];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[125] = chanx_right_in[124];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[126] = chanx_right_in[125];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[127] = chanx_right_in[126];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[129] = chanx_right_in[128];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[130] = chanx_right_in[129];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[131] = chanx_right_in[130];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[133] = chanx_right_in[132];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[134] = chanx_right_in[133];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[135] = chanx_right_in[134];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[137] = chanx_right_in[136];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[138] = chanx_right_in[137];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[139] = chanx_right_in[138];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[141] = chanx_right_in[140];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[142] = chanx_right_in[141];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[143] = chanx_right_in[142];
// ----- Local connection due to Wire 330 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[145] = chanx_right_in[144];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[146] = chanx_right_in[145];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[147] = chanx_right_in[146];
// ----- Local connection due to Wire 334 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[149] = chanx_right_in[148];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[1];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[5];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[9];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 419 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 420 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 423 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 424 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 428 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 432 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 436 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[83] = chanx_left_in[82];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 440 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[87] = chanx_left_in[86];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[91] = chanx_left_in[90];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- Local connection due to Wire 448 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[95] = chanx_left_in[94];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[97] = chanx_left_in[96];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[98] = chanx_left_in[97];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[99] = chanx_left_in[98];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[101] = chanx_left_in[100];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[102] = chanx_left_in[101];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[103] = chanx_left_in[102];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[105] = chanx_left_in[104];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[106] = chanx_left_in[105];
// ----- Local connection due to Wire 460 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[107] = chanx_left_in[106];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[109] = chanx_left_in[108];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[110] = chanx_left_in[109];
// ----- Local connection due to Wire 464 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[111] = chanx_left_in[110];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[113] = chanx_left_in[112];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[114] = chanx_left_in[113];
// ----- Local connection due to Wire 468 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[115] = chanx_left_in[114];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[117] = chanx_left_in[116];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[118] = chanx_left_in[117];
// ----- Local connection due to Wire 472 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[119] = chanx_left_in[118];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[121] = chanx_left_in[120];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[122] = chanx_left_in[121];
// ----- Local connection due to Wire 476 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[123] = chanx_left_in[122];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[125] = chanx_left_in[124];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[126] = chanx_left_in[125];
// ----- Local connection due to Wire 480 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[127] = chanx_left_in[126];
// ----- Local connection due to Wire 482 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[129] = chanx_left_in[128];
// ----- Local connection due to Wire 483 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[130] = chanx_left_in[129];
// ----- Local connection due to Wire 484 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[131] = chanx_left_in[130];
// ----- Local connection due to Wire 486 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[133] = chanx_left_in[132];
// ----- Local connection due to Wire 487 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[134] = chanx_left_in[133];
// ----- Local connection due to Wire 488 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[135] = chanx_left_in[134];
// ----- Local connection due to Wire 490 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[137] = chanx_left_in[136];
// ----- Local connection due to Wire 491 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[138] = chanx_left_in[137];
// ----- Local connection due to Wire 492 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[139] = chanx_left_in[138];
// ----- Local connection due to Wire 494 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[141] = chanx_left_in[140];
// ----- Local connection due to Wire 495 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[142] = chanx_left_in[141];
// ----- Local connection due to Wire 496 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[143] = chanx_left_in[142];
// ----- Local connection due to Wire 498 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[145] = chanx_left_in[144];
// ----- Local connection due to Wire 499 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[146] = chanx_left_in[145];
// ----- Local connection due to Wire 500 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[147] = chanx_left_in[146];
// ----- Local connection due to Wire 502 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[149] = chanx_left_in[148];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size8 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[1], chanx_right_in[7], chanx_left_in[0], chanx_left_in[3]}),
		.sram(mux_2level_tapbuf_size8_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_0_sram_inv[0:5]),
		.out(chany_top_out[0]));

	mux_2level_tapbuf_size8 mux_right_track_288 (
		.in({chany_top_in[35], chany_top_in[73], chany_top_in[111], chany_top_in[149], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[48], chanx_left_in[98]}),
		.sram(mux_2level_tapbuf_size8_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_1_sram_inv[0:5]),
		.out(chanx_right_out[144]));

	mux_2level_tapbuf_size8 mux_left_track_9 (
		.in({chany_top_in[37], chany_top_in[75], chany_top_in[113], chanx_right_in[1], chanx_right_in[52], chanx_right_in[102], left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_2_sram_inv[0:5]),
		.out(chanx_left_out[4]));

	mux_2level_tapbuf_size8 mux_left_track_17 (
		.in({chany_top_in[36], chany_top_in[74], chany_top_in[112], chanx_right_in[2], chanx_right_in[53], chanx_right_in[104], left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_3_sram_inv[0:5]),
		.out(chanx_left_out[8]));

	mux_2level_tapbuf_size8 mux_left_track_49 (
		.in({chany_top_in[32], chany_top_in[70], chany_top_in[108], chany_top_in[146], chanx_right_in[8], chanx_right_in[58], chanx_right_in[109], left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_4_sram_inv[0:5]),
		.out(chanx_left_out[24]));

	mux_2level_tapbuf_size8 mux_left_track_57 (
		.in({chany_top_in[31], chany_top_in[69], chany_top_in[107], chany_top_in[145], chanx_right_in[9], chanx_right_in[60], chanx_right_in[110], left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_5_sram_inv[0:5]),
		.out(chanx_left_out[28]));

	mux_2level_tapbuf_size8 mux_left_track_73 (
		.in({chany_top_in[29], chany_top_in[67], chany_top_in[105], chany_top_in[143], chanx_right_in[12], chanx_right_in[62], chanx_right_in[113], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_6_sram_inv[0:5]),
		.out(chanx_left_out[36]));

	mux_2level_tapbuf_size8 mux_left_track_81 (
		.in({chany_top_in[28], chany_top_in[66], chany_top_in[104], chany_top_in[142], chanx_right_in[13], chanx_right_in[64], chanx_right_in[114], left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_7_sram_inv[0:5]),
		.out(chanx_left_out[40]));

	mux_2level_tapbuf_size8 mux_left_track_89 (
		.in({chany_top_in[27], chany_top_in[65], chany_top_in[103], chany_top_in[141], chanx_right_in[14], chanx_right_in[65], chanx_right_in[116], left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_8_sram_inv[0:5]),
		.out(chanx_left_out[44]));

	mux_2level_tapbuf_size8 mux_left_track_97 (
		.in({chany_top_in[26], chany_top_in[64], chany_top_in[102], chany_top_in[140], chanx_right_in[16], chanx_right_in[66], chanx_right_in[117], left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_9_sram_inv[0:5]),
		.out(chanx_left_out[48]));

	mux_2level_tapbuf_size8 mux_left_track_105 (
		.in({chany_top_in[25], chany_top_in[63], chany_top_in[101], chany_top_in[139], chanx_right_in[17], chanx_right_in[68], chanx_right_in[118], left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_10_sram_inv[0:5]),
		.out(chanx_left_out[52]));

	mux_2level_tapbuf_size8 mux_left_track_113 (
		.in({chany_top_in[24], chany_top_in[62], chany_top_in[100], chany_top_in[138], chanx_right_in[18], chanx_right_in[69], chanx_right_in[120], left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_11_sram_inv[0:5]),
		.out(chanx_left_out[56]));

	mux_2level_tapbuf_size8 mux_left_track_121 (
		.in({chany_top_in[23], chany_top_in[61], chany_top_in[99], chany_top_in[137], chanx_right_in[20], chanx_right_in[70], chanx_right_in[121], left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_12_sram_inv[0:5]),
		.out(chanx_left_out[60]));

	mux_2level_tapbuf_size8 mux_left_track_129 (
		.in({chany_top_in[22], chany_top_in[60], chany_top_in[98], chany_top_in[136], chanx_right_in[21], chanx_right_in[72], chanx_right_in[122], left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_13_sram_inv[0:5]),
		.out(chanx_left_out[64]));

	mux_2level_tapbuf_size8 mux_left_track_145 (
		.in({chany_top_in[20], chany_top_in[58], chany_top_in[96], chany_top_in[134], chanx_right_in[24], chanx_right_in[74], chanx_right_in[125], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_14_sram_inv[0:5]),
		.out(chanx_left_out[72]));

	mux_2level_tapbuf_size8 mux_left_track_153 (
		.in({chany_top_in[19], chany_top_in[57], chany_top_in[95], chany_top_in[133], chanx_right_in[25], chanx_right_in[76], chanx_right_in[126], left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_15_sram_inv[0:5]),
		.out(chanx_left_out[76]));

	mux_2level_tapbuf_size8 mux_left_track_161 (
		.in({chany_top_in[18], chany_top_in[56], chany_top_in[94], chany_top_in[132], chanx_right_in[26], chanx_right_in[77], chanx_right_in[128], left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_16_sram_inv[0:5]),
		.out(chanx_left_out[80]));

	mux_2level_tapbuf_size8 mux_left_track_169 (
		.in({chany_top_in[17], chany_top_in[55], chany_top_in[93], chany_top_in[131], chanx_right_in[28], chanx_right_in[78], chanx_right_in[129], left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_17_sram_inv[0:5]),
		.out(chanx_left_out[84]));

	mux_2level_tapbuf_size8 mux_left_track_177 (
		.in({chany_top_in[16], chany_top_in[54], chany_top_in[92], chany_top_in[130], chanx_right_in[29], chanx_right_in[80], chanx_right_in[130], left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_18_sram_inv[0:5]),
		.out(chanx_left_out[88]));

	mux_2level_tapbuf_size8 mux_left_track_185 (
		.in({chany_top_in[15], chany_top_in[53], chany_top_in[91], chany_top_in[129], chanx_right_in[30], chanx_right_in[81], chanx_right_in[132], left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_19_sram_inv[0:5]),
		.out(chanx_left_out[92]));

	mux_2level_tapbuf_size8 mux_left_track_193 (
		.in({chany_top_in[14], chany_top_in[52], chany_top_in[90], chany_top_in[128], chanx_right_in[32], chanx_right_in[82], chanx_right_in[133], left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_20_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_20_sram_inv[0:5]),
		.out(chanx_left_out[96]));

	mux_2level_tapbuf_size8 mux_left_track_201 (
		.in({chany_top_in[13], chany_top_in[51], chany_top_in[89], chany_top_in[127], chanx_right_in[33], chanx_right_in[84], chanx_right_in[134], left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_21_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_21_sram_inv[0:5]),
		.out(chanx_left_out[100]));

	mux_2level_tapbuf_size8 mux_left_track_217 (
		.in({chany_top_in[11], chany_top_in[49], chany_top_in[87], chany_top_in[125], chanx_right_in[36], chanx_right_in[86], chanx_right_in[137], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_22_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_22_sram_inv[0:5]),
		.out(chanx_left_out[108]));

	mux_2level_tapbuf_size8 mux_left_track_225 (
		.in({chany_top_in[10], chany_top_in[48], chany_top_in[86], chany_top_in[124], chanx_right_in[37], chanx_right_in[88], chanx_right_in[138], left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_23_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_23_sram_inv[0:5]),
		.out(chanx_left_out[112]));

	mux_2level_tapbuf_size8 mux_left_track_233 (
		.in({chany_top_in[9], chany_top_in[47], chany_top_in[85], chany_top_in[123], chanx_right_in[38], chanx_right_in[89], chanx_right_in[140], left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_24_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_24_sram_inv[0:5]),
		.out(chanx_left_out[116]));

	mux_2level_tapbuf_size8 mux_left_track_241 (
		.in({chany_top_in[8], chany_top_in[46], chany_top_in[84], chany_top_in[122], chanx_right_in[40], chanx_right_in[90], chanx_right_in[141], left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_25_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_25_sram_inv[0:5]),
		.out(chanx_left_out[120]));

	mux_2level_tapbuf_size8 mux_left_track_249 (
		.in({chany_top_in[7], chany_top_in[45], chany_top_in[83], chany_top_in[121], chanx_right_in[41], chanx_right_in[92], chanx_right_in[142], left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_26_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_26_sram_inv[0:5]),
		.out(chanx_left_out[124]));

	mux_2level_tapbuf_size8 mux_left_track_257 (
		.in({chany_top_in[6], chany_top_in[44], chany_top_in[82], chany_top_in[120], chanx_right_in[42], chanx_right_in[93], chanx_right_in[144], left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_27_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_27_sram_inv[0:5]),
		.out(chanx_left_out[128]));

	mux_2level_tapbuf_size8 mux_left_track_265 (
		.in({chany_top_in[5], chany_top_in[43], chany_top_in[81], chany_top_in[119], chanx_right_in[44], chanx_right_in[94], chanx_right_in[145], left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_28_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_28_sram_inv[0:5]),
		.out(chanx_left_out[132]));

	mux_2level_tapbuf_size8 mux_left_track_273 (
		.in({chany_top_in[4], chany_top_in[42], chany_top_in[80], chany_top_in[118], chanx_right_in[45], chanx_right_in[96], chanx_right_in[146], left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_29_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_29_sram_inv[0:5]),
		.out(chanx_left_out[136]));

	mux_2level_tapbuf_size8_mem mem_top_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_0_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_1_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_2_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_3_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_4_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_5_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_6_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_7_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_8_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_97 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_9_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_105 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_10_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_113 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_11_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_121 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_12_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_129 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_13_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_145 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_14_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_153 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_15_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_161 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_16_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_169 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_17_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_177 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_18_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_185 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_19_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_193 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_20_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_20_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_201 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_21_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_21_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_217 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_22_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_22_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_225 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_23_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_23_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_233 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_24_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_24_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_241 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_25_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_25_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_249 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_26_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_26_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_257 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_27_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_27_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_265 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_28_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_28_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_273 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_29_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_29_sram_inv[0:5]));

	mux_2level_tapbuf_size6 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_right_in[2], chanx_right_in[11]}),
		.sram(mux_2level_tapbuf_size6_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_0_sram_inv[0:5]),
		.out(chany_top_out[1]));

	mux_2level_tapbuf_size6 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_right_in[4], chanx_right_in[15]}),
		.sram(mux_2level_tapbuf_size6_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_1_sram_inv[0:5]),
		.out(chany_top_out[2]));

	mux_2level_tapbuf_size6 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_right_in[5], chanx_right_in[19]}),
		.sram(mux_2level_tapbuf_size6_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_2_sram_inv[0:5]),
		.out(chany_top_out[3]));

	mux_2level_tapbuf_size6 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_right_in[6], chanx_right_in[23]}),
		.sram(mux_2level_tapbuf_size6_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_3_sram_inv[0:5]),
		.out(chany_top_out[4]));

	mux_2level_tapbuf_size6 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_right_in[8], chanx_right_in[27]}),
		.sram(mux_2level_tapbuf_size6_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_4_sram_inv[0:5]),
		.out(chany_top_out[5]));

	mux_2level_tapbuf_size6 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[14], chanx_right_in[47]}),
		.sram(mux_2level_tapbuf_size6_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_5_sram_inv[0:5]),
		.out(chany_top_out[10]));

	mux_2level_tapbuf_size6 mux_top_track_22 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_right_in[16], chanx_right_in[51]}),
		.sram(mux_2level_tapbuf_size6_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_6_sram_inv[0:5]),
		.out(chany_top_out[11]));

	mux_2level_tapbuf_size6 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_right_in[17], chanx_right_in[55]}),
		.sram(mux_2level_tapbuf_size6_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_7_sram_inv[0:5]),
		.out(chany_top_out[12]));

	mux_2level_tapbuf_size6 mux_top_track_26 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_right_in[18], chanx_right_in[59]}),
		.sram(mux_2level_tapbuf_size6_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_8_sram_inv[0:5]),
		.out(chany_top_out[13]));

	mux_2level_tapbuf_size6 mux_top_track_28 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_right_in[20], chanx_right_in[63]}),
		.sram(mux_2level_tapbuf_size6_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_9_sram_inv[0:5]),
		.out(chany_top_out[14]));

	mux_2level_tapbuf_size6 mux_top_track_30 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_right_in[21], chanx_right_in[67]}),
		.sram(mux_2level_tapbuf_size6_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_10_sram_inv[0:5]),
		.out(chany_top_out[15]));

	mux_2level_tapbuf_size6 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[28], chanx_right_in[87]}),
		.sram(mux_2level_tapbuf_size6_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_11_sram_inv[0:5]),
		.out(chany_top_out[20]));

	mux_2level_tapbuf_size6 mux_top_track_42 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_right_in[29], chanx_right_in[91]}),
		.sram(mux_2level_tapbuf_size6_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_12_sram_inv[0:5]),
		.out(chany_top_out[21]));

	mux_2level_tapbuf_size6 mux_top_track_44 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_right_in[30], chanx_right_in[95]}),
		.sram(mux_2level_tapbuf_size6_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_13_sram_inv[0:5]),
		.out(chany_top_out[22]));

	mux_2level_tapbuf_size6 mux_top_track_46 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_right_in[32], chanx_right_in[99]}),
		.sram(mux_2level_tapbuf_size6_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_14_sram_inv[0:5]),
		.out(chany_top_out[23]));

	mux_2level_tapbuf_size6 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_right_in[33], chanx_right_in[103]}),
		.sram(mux_2level_tapbuf_size6_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_15_sram_inv[0:5]),
		.out(chany_top_out[24]));

	mux_2level_tapbuf_size6 mux_top_track_50 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_right_in[34], chanx_right_in[107]}),
		.sram(mux_2level_tapbuf_size6_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_16_sram_inv[0:5]),
		.out(chany_top_out[25]));

	mux_2level_tapbuf_size6 mux_top_track_60 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[41], chanx_right_in[127]}),
		.sram(mux_2level_tapbuf_size6_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_17_sram_inv[0:5]),
		.out(chany_top_out[30]));

	mux_2level_tapbuf_size6 mux_top_track_62 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_right_in[42], chanx_right_in[131]}),
		.sram(mux_2level_tapbuf_size6_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_18_sram_inv[0:5]),
		.out(chany_top_out[31]));

	mux_2level_tapbuf_size6 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_right_in[44], chanx_right_in[135]}),
		.sram(mux_2level_tapbuf_size6_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_19_sram_inv[0:5]),
		.out(chany_top_out[32]));

	mux_2level_tapbuf_size6 mux_top_track_66 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_right_in[45], chanx_right_in[139]}),
		.sram(mux_2level_tapbuf_size6_20_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_20_sram_inv[0:5]),
		.out(chany_top_out[33]));

	mux_2level_tapbuf_size6 mux_top_track_68 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_right_in[46], chanx_right_in[143]}),
		.sram(mux_2level_tapbuf_size6_21_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_21_sram_inv[0:5]),
		.out(chany_top_out[34]));

	mux_2level_tapbuf_size6 mux_top_track_70 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_right_in[48], chanx_right_in[147]}),
		.sram(mux_2level_tapbuf_size6_22_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_22_sram_inv[0:5]),
		.out(chany_top_out[35]));

	mux_2level_tapbuf_size6 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[54], chanx_left_in[146]}),
		.sram(mux_2level_tapbuf_size6_23_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_23_sram_inv[0:5]),
		.out(chany_top_out[40]));

	mux_2level_tapbuf_size6 mux_top_track_82 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_right_in[56], chanx_left_in[145]}),
		.sram(mux_2level_tapbuf_size6_24_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_24_sram_inv[0:5]),
		.out(chany_top_out[41]));

	mux_2level_tapbuf_size6 mux_top_track_84 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_right_in[57], chanx_left_in[144]}),
		.sram(mux_2level_tapbuf_size6_25_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_25_sram_inv[0:5]),
		.out(chany_top_out[42]));

	mux_2level_tapbuf_size6 mux_top_track_86 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_right_in[58], chanx_left_in[142]}),
		.sram(mux_2level_tapbuf_size6_26_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_26_sram_inv[0:5]),
		.out(chany_top_out[43]));

	mux_2level_tapbuf_size6 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_right_in[60], chanx_left_in[141]}),
		.sram(mux_2level_tapbuf_size6_27_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_27_sram_inv[0:5]),
		.out(chany_top_out[44]));

	mux_2level_tapbuf_size6 mux_top_track_90 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_right_in[61], chanx_left_in[140]}),
		.sram(mux_2level_tapbuf_size6_28_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_28_sram_inv[0:5]),
		.out(chany_top_out[45]));

	mux_2level_tapbuf_size6 mux_top_track_100 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[68], chanx_left_in[133]}),
		.sram(mux_2level_tapbuf_size6_29_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_29_sram_inv[0:5]),
		.out(chany_top_out[50]));

	mux_2level_tapbuf_size6 mux_top_track_102 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_right_in[69], chanx_left_in[132]}),
		.sram(mux_2level_tapbuf_size6_30_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_30_sram_inv[0:5]),
		.out(chany_top_out[51]));

	mux_2level_tapbuf_size6 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_right_in[70], chanx_left_in[130]}),
		.sram(mux_2level_tapbuf_size6_31_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_31_sram_inv[0:5]),
		.out(chany_top_out[52]));

	mux_2level_tapbuf_size6 mux_top_track_106 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_right_in[72], chanx_left_in[129]}),
		.sram(mux_2level_tapbuf_size6_32_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_32_sram_inv[0:5]),
		.out(chany_top_out[53]));

	mux_2level_tapbuf_size6 mux_top_track_108 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_right_in[73], chanx_left_in[128]}),
		.sram(mux_2level_tapbuf_size6_33_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_33_sram_inv[0:5]),
		.out(chany_top_out[54]));

	mux_2level_tapbuf_size6 mux_top_track_110 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_right_in[74], chanx_left_in[126]}),
		.sram(mux_2level_tapbuf_size6_34_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_34_sram_inv[0:5]),
		.out(chany_top_out[55]));

	mux_2level_tapbuf_size6 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[81], chanx_left_in[120]}),
		.sram(mux_2level_tapbuf_size6_35_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_35_sram_inv[0:5]),
		.out(chany_top_out[60]));

	mux_2level_tapbuf_size6 mux_top_track_122 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_right_in[82], chanx_left_in[118]}),
		.sram(mux_2level_tapbuf_size6_36_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_36_sram_inv[0:5]),
		.out(chany_top_out[61]));

	mux_2level_tapbuf_size6 mux_top_track_124 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_right_in[84], chanx_left_in[117]}),
		.sram(mux_2level_tapbuf_size6_37_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_37_sram_inv[0:5]),
		.out(chany_top_out[62]));

	mux_2level_tapbuf_size6 mux_top_track_126 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_right_in[85], chanx_left_in[116]}),
		.sram(mux_2level_tapbuf_size6_38_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_38_sram_inv[0:5]),
		.out(chany_top_out[63]));

	mux_2level_tapbuf_size6 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_right_in[86], chanx_left_in[114]}),
		.sram(mux_2level_tapbuf_size6_39_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_39_sram_inv[0:5]),
		.out(chany_top_out[64]));

	mux_2level_tapbuf_size6 mux_top_track_130 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_right_in[88], chanx_left_in[113]}),
		.sram(mux_2level_tapbuf_size6_40_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_40_sram_inv[0:5]),
		.out(chany_top_out[65]));

	mux_2level_tapbuf_size6 mux_top_track_140 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[94], chanx_left_in[106]}),
		.sram(mux_2level_tapbuf_size6_41_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_41_sram_inv[0:5]),
		.out(chany_top_out[70]));

	mux_2level_tapbuf_size6 mux_top_track_142 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_right_in[96], chanx_left_in[105]}),
		.sram(mux_2level_tapbuf_size6_42_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_42_sram_inv[0:5]),
		.out(chany_top_out[71]));

	mux_2level_tapbuf_size6 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_right_in[97], chanx_left_in[104]}),
		.sram(mux_2level_tapbuf_size6_43_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_43_sram_inv[0:5]),
		.out(chany_top_out[72]));

	mux_2level_tapbuf_size6 mux_top_track_146 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_right_in[98], chanx_left_in[102]}),
		.sram(mux_2level_tapbuf_size6_44_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_44_sram_inv[0:5]),
		.out(chany_top_out[73]));

	mux_2level_tapbuf_size6 mux_top_track_148 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_right_in[100], chanx_left_in[101]}),
		.sram(mux_2level_tapbuf_size6_45_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_45_sram_inv[0:5]),
		.out(chany_top_out[74]));

	mux_2level_tapbuf_size6 mux_top_track_150 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_right_in[101], chanx_left_in[100]}),
		.sram(mux_2level_tapbuf_size6_46_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_46_sram_inv[0:5]),
		.out(chany_top_out[75]));

	mux_2level_tapbuf_size6 mux_top_track_160 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[108], chanx_left_in[93]}),
		.sram(mux_2level_tapbuf_size6_47_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_47_sram_inv[0:5]),
		.out(chany_top_out[80]));

	mux_2level_tapbuf_size6 mux_top_track_162 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_right_in[109], chanx_left_in[92]}),
		.sram(mux_2level_tapbuf_size6_48_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_48_sram_inv[0:5]),
		.out(chany_top_out[81]));

	mux_2level_tapbuf_size6 mux_top_track_164 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_right_in[110], chanx_left_in[90]}),
		.sram(mux_2level_tapbuf_size6_49_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_49_sram_inv[0:5]),
		.out(chany_top_out[82]));

	mux_2level_tapbuf_size6 mux_top_track_166 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_right_in[112], chanx_left_in[89]}),
		.sram(mux_2level_tapbuf_size6_50_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_50_sram_inv[0:5]),
		.out(chany_top_out[83]));

	mux_2level_tapbuf_size6 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_right_in[113], chanx_left_in[88]}),
		.sram(mux_2level_tapbuf_size6_51_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_51_sram_inv[0:5]),
		.out(chany_top_out[84]));

	mux_2level_tapbuf_size6 mux_top_track_170 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_right_in[114], chanx_left_in[86]}),
		.sram(mux_2level_tapbuf_size6_52_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_52_sram_inv[0:5]),
		.out(chany_top_out[85]));

	mux_2level_tapbuf_size6 mux_top_track_180 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[121], chanx_left_in[80]}),
		.sram(mux_2level_tapbuf_size6_53_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_53_sram_inv[0:5]),
		.out(chany_top_out[90]));

	mux_2level_tapbuf_size6 mux_top_track_182 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_right_in[122], chanx_left_in[78]}),
		.sram(mux_2level_tapbuf_size6_54_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_54_sram_inv[0:5]),
		.out(chany_top_out[91]));

	mux_2level_tapbuf_size6 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_right_in[124], chanx_left_in[77]}),
		.sram(mux_2level_tapbuf_size6_55_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_55_sram_inv[0:5]),
		.out(chany_top_out[92]));

	mux_2level_tapbuf_size6 mux_top_track_186 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_right_in[125], chanx_left_in[76]}),
		.sram(mux_2level_tapbuf_size6_56_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_56_sram_inv[0:5]),
		.out(chany_top_out[93]));

	mux_2level_tapbuf_size6 mux_top_track_188 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_right_in[126], chanx_left_in[74]}),
		.sram(mux_2level_tapbuf_size6_57_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_57_sram_inv[0:5]),
		.out(chany_top_out[94]));

	mux_2level_tapbuf_size6 mux_top_track_190 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_right_in[128], chanx_left_in[73]}),
		.sram(mux_2level_tapbuf_size6_58_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_58_sram_inv[0:5]),
		.out(chany_top_out[95]));

	mux_2level_tapbuf_size6 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[134], chanx_left_in[66]}),
		.sram(mux_2level_tapbuf_size6_59_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_59_sram_inv[0:5]),
		.out(chany_top_out[100]));

	mux_2level_tapbuf_size6 mux_top_track_202 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_right_in[136], chanx_left_in[65]}),
		.sram(mux_2level_tapbuf_size6_60_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_60_sram_inv[0:5]),
		.out(chany_top_out[101]));

	mux_2level_tapbuf_size6 mux_top_track_204 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_right_in[137], chanx_left_in[64]}),
		.sram(mux_2level_tapbuf_size6_61_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_61_sram_inv[0:5]),
		.out(chany_top_out[102]));

	mux_2level_tapbuf_size6 mux_top_track_206 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_right_in[138], chanx_left_in[62]}),
		.sram(mux_2level_tapbuf_size6_62_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_62_sram_inv[0:5]),
		.out(chany_top_out[103]));

	mux_2level_tapbuf_size6 mux_top_track_208 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_right_in[140], chanx_left_in[61]}),
		.sram(mux_2level_tapbuf_size6_63_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_63_sram_inv[0:5]),
		.out(chany_top_out[104]));

	mux_2level_tapbuf_size6 mux_top_track_210 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_right_in[141], chanx_left_in[60]}),
		.sram(mux_2level_tapbuf_size6_64_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_64_sram_inv[0:5]),
		.out(chany_top_out[105]));

	mux_2level_tapbuf_size6 mux_top_track_220 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_right_in[148], chanx_left_in[53]}),
		.sram(mux_2level_tapbuf_size6_65_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_65_sram_inv[0:5]),
		.out(chany_top_out[110]));

	mux_2level_tapbuf_size6 mux_top_track_226 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_left_in[49], chanx_left_in[149]}),
		.sram(mux_2level_tapbuf_size6_66_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_66_sram_inv[0:5]),
		.out(chany_top_out[113]));

	mux_2level_tapbuf_size6 mux_top_track_228 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_left_in[48], chanx_left_in[147]}),
		.sram(mux_2level_tapbuf_size6_67_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_67_sram_inv[0:5]),
		.out(chany_top_out[114]));

	mux_2level_tapbuf_size6 mux_top_track_230 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_left_in[46], chanx_left_in[143]}),
		.sram(mux_2level_tapbuf_size6_68_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_68_sram_inv[0:5]),
		.out(chany_top_out[115]));

	mux_2level_tapbuf_size6 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_left_in[40], chanx_left_in[123]}),
		.sram(mux_2level_tapbuf_size6_69_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_69_sram_inv[0:5]),
		.out(chany_top_out[120]));

	mux_2level_tapbuf_size6 mux_top_track_242 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_left_in[38], chanx_left_in[119]}),
		.sram(mux_2level_tapbuf_size6_70_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_70_sram_inv[0:5]),
		.out(chany_top_out[121]));

	mux_2level_tapbuf_size6 mux_top_track_244 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_left_in[37], chanx_left_in[115]}),
		.sram(mux_2level_tapbuf_size6_71_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_71_sram_inv[0:5]),
		.out(chany_top_out[122]));

	mux_2level_tapbuf_size6 mux_top_track_246 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_left_in[36], chanx_left_in[111]}),
		.sram(mux_2level_tapbuf_size6_72_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_72_sram_inv[0:5]),
		.out(chany_top_out[123]));

	mux_2level_tapbuf_size6 mux_top_track_248 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_left_in[34], chanx_left_in[107]}),
		.sram(mux_2level_tapbuf_size6_73_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_73_sram_inv[0:5]),
		.out(chany_top_out[124]));

	mux_2level_tapbuf_size6 mux_top_track_250 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_left_in[33], chanx_left_in[103]}),
		.sram(mux_2level_tapbuf_size6_74_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_74_sram_inv[0:5]),
		.out(chany_top_out[125]));

	mux_2level_tapbuf_size6 mux_top_track_260 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_left_in[26], chanx_left_in[83]}),
		.sram(mux_2level_tapbuf_size6_75_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_75_sram_inv[0:5]),
		.out(chany_top_out[130]));

	mux_2level_tapbuf_size6 mux_top_track_262 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_left_in[25], chanx_left_in[79]}),
		.sram(mux_2level_tapbuf_size6_76_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_76_sram_inv[0:5]),
		.out(chany_top_out[131]));

	mux_2level_tapbuf_size6 mux_top_track_264 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_left_in[24], chanx_left_in[75]}),
		.sram(mux_2level_tapbuf_size6_77_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_77_sram_inv[0:5]),
		.out(chany_top_out[132]));

	mux_2level_tapbuf_size6 mux_top_track_266 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_left_in[22], chanx_left_in[71]}),
		.sram(mux_2level_tapbuf_size6_78_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_78_sram_inv[0:5]),
		.out(chany_top_out[133]));

	mux_2level_tapbuf_size6 mux_top_track_268 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_left_in[21], chanx_left_in[67]}),
		.sram(mux_2level_tapbuf_size6_79_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_79_sram_inv[0:5]),
		.out(chany_top_out[134]));

	mux_2level_tapbuf_size6 mux_top_track_270 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_left_in[20], chanx_left_in[63]}),
		.sram(mux_2level_tapbuf_size6_80_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_80_sram_inv[0:5]),
		.out(chany_top_out[135]));

	mux_2level_tapbuf_size6 mux_top_track_280 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_30_, chanx_left_in[13], chanx_left_in[43]}),
		.sram(mux_2level_tapbuf_size6_81_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_81_sram_inv[0:5]),
		.out(chany_top_out[140]));

	mux_2level_tapbuf_size6 mux_top_track_282 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_left_in[12], chanx_left_in[39]}),
		.sram(mux_2level_tapbuf_size6_82_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_82_sram_inv[0:5]),
		.out(chany_top_out[141]));

	mux_2level_tapbuf_size6 mux_top_track_284 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_left_in[10], chanx_left_in[35]}),
		.sram(mux_2level_tapbuf_size6_83_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_83_sram_inv[0:5]),
		.out(chany_top_out[142]));

	mux_2level_tapbuf_size6 mux_top_track_286 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_33_, chanx_left_in[9], chanx_left_in[31]}),
		.sram(mux_2level_tapbuf_size6_84_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_84_sram_inv[0:5]),
		.out(chany_top_out[143]));

	mux_2level_tapbuf_size6 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_34_, chanx_left_in[8], chanx_left_in[27]}),
		.sram(mux_2level_tapbuf_size6_85_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_85_sram_inv[0:5]),
		.out(chany_top_out[144]));

	mux_2level_tapbuf_size6 mux_top_track_290 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_35_, chanx_left_in[6], chanx_left_in[23]}),
		.sram(mux_2level_tapbuf_size6_86_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_86_sram_inv[0:5]),
		.out(chany_top_out[145]));

	mux_2level_tapbuf_size6_mem mem_top_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_0_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_1_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_6 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_2_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_3_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_4_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_5_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_22 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_6_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_7_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_8_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_9_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_30 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_10_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_11_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_12_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_13_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_46 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_14_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_15_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_16_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_17_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_62 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_18_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_19_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_20_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_20_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_21_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_21_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_70 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_22_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_22_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_23_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_23_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_24_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_24_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_25_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_25_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_86 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_26_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_26_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_27_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_27_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_28_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_28_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_29_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_29_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_102 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_30_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_30_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_31_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_31_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_106 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_32_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_32_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_33_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_33_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_110 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_34_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_34_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_35_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_35_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_36_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_36_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_124 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_37_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_37_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_126 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_38_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_38_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_39_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_39_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_40_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_40_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_41_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_41_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_142 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_42_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_42_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_43_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_43_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_44_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_44_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_45_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_45_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_150 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_46_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_46_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_47_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_47_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_48_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_48_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_49_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_49_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_166 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_50_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_50_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_51_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_51_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_52_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_52_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_53_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_53_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_182 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_54_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_54_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_55_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_55_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_56_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_56_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_57_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_57_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_190 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_58_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_58_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_59_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_59_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_60_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_60_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_61_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_61_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_206 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_62_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_62_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_63_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_63_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_210 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_64_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_64_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_220 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_65_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_65_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_226 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_66_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_66_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_228 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_67_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_67_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_230 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_68_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_68_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_69_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_69_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_242 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_70_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_70_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_244 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_71_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_71_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_246 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_72_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_72_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_73_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_73_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_250 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_74_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_74_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_260 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_75_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_75_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_262 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_76_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_76_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_77_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_77_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_266 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_78_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_78_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_268 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_78_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_79_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_79_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_79_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_270 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_79_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_80_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_80_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_80_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_81_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_81_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_81_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_282 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_81_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_82_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_82_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_82_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_284 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_82_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_83_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_83_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_83_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_286 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_83_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_84_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_84_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_84_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_84_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_85_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_85_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_85_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_290 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_85_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_86_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_86_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_86_sram_inv[0:5]));

	mux_2level_tapbuf_size5 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_right_in[9], chanx_right_in[31]}),
		.sram(mux_2level_tapbuf_size5_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_0_sram_inv[0:5]),
		.out(chany_top_out[6]));

	mux_2level_tapbuf_size5 mux_top_track_14 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_right_in[10], chanx_right_in[35]}),
		.sram(mux_2level_tapbuf_size5_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_1_sram_inv[0:5]),
		.out(chany_top_out[7]));

	mux_2level_tapbuf_size5 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_right_in[12], chanx_right_in[39]}),
		.sram(mux_2level_tapbuf_size5_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_2_sram_inv[0:5]),
		.out(chany_top_out[8]));

	mux_2level_tapbuf_size5 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[13], chanx_right_in[43]}),
		.sram(mux_2level_tapbuf_size5_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_3_sram_inv[0:5]),
		.out(chany_top_out[9]));

	mux_2level_tapbuf_size5 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_right_in[22], chanx_right_in[71]}),
		.sram(mux_2level_tapbuf_size5_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_4_sram_inv[0:5]),
		.out(chany_top_out[16]));

	mux_2level_tapbuf_size5 mux_top_track_34 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_right_in[24], chanx_right_in[75]}),
		.sram(mux_2level_tapbuf_size5_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_5_sram_inv[0:5]),
		.out(chany_top_out[17]));

	mux_2level_tapbuf_size5 mux_top_track_36 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_right_in[25], chanx_right_in[79]}),
		.sram(mux_2level_tapbuf_size5_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_6_sram_inv[0:5]),
		.out(chany_top_out[18]));

	mux_2level_tapbuf_size5 mux_top_track_38 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[26], chanx_right_in[83]}),
		.sram(mux_2level_tapbuf_size5_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_7_sram_inv[0:5]),
		.out(chany_top_out[19]));

	mux_2level_tapbuf_size5 mux_top_track_52 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_right_in[36], chanx_right_in[111]}),
		.sram(mux_2level_tapbuf_size5_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_8_sram_inv[0:5]),
		.out(chany_top_out[26]));

	mux_2level_tapbuf_size5 mux_top_track_54 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_right_in[37], chanx_right_in[115]}),
		.sram(mux_2level_tapbuf_size5_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_9_sram_inv[0:5]),
		.out(chany_top_out[27]));

	mux_2level_tapbuf_size5 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_right_in[38], chanx_right_in[119]}),
		.sram(mux_2level_tapbuf_size5_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_10_sram_inv[0:5]),
		.out(chany_top_out[28]));

	mux_2level_tapbuf_size5 mux_top_track_58 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[40], chanx_right_in[123]}),
		.sram(mux_2level_tapbuf_size5_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_11_sram_inv[0:5]),
		.out(chany_top_out[29]));

	mux_2level_tapbuf_size5 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_right_in[49], chanx_right_in[149]}),
		.sram(mux_2level_tapbuf_size5_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_12_sram_inv[0:5]),
		.out(chany_top_out[36]));

	mux_2level_tapbuf_size5 mux_top_track_78 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[53], chanx_left_in[148]}),
		.sram(mux_2level_tapbuf_size5_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_13_sram_inv[0:5]),
		.out(chany_top_out[39]));

	mux_2level_tapbuf_size5 mux_top_track_92 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_right_in[62], chanx_left_in[138]}),
		.sram(mux_2level_tapbuf_size5_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_14_sram_inv[0:5]),
		.out(chany_top_out[46]));

	mux_2level_tapbuf_size5 mux_top_track_94 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_right_in[64], chanx_left_in[137]}),
		.sram(mux_2level_tapbuf_size5_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_15_sram_inv[0:5]),
		.out(chany_top_out[47]));

	mux_2level_tapbuf_size5 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_right_in[65], chanx_left_in[136]}),
		.sram(mux_2level_tapbuf_size5_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_16_sram_inv[0:5]),
		.out(chany_top_out[48]));

	mux_2level_tapbuf_size5 mux_top_track_98 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[66], chanx_left_in[134]}),
		.sram(mux_2level_tapbuf_size5_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_17_sram_inv[0:5]),
		.out(chany_top_out[49]));

	mux_2level_tapbuf_size5 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_right_in[76], chanx_left_in[125]}),
		.sram(mux_2level_tapbuf_size5_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_18_sram_inv[0:5]),
		.out(chany_top_out[56]));

	mux_2level_tapbuf_size5 mux_top_track_114 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_right_in[77], chanx_left_in[124]}),
		.sram(mux_2level_tapbuf_size5_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_19_sram_inv[0:5]),
		.out(chany_top_out[57]));

	mux_2level_tapbuf_size5 mux_top_track_116 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_right_in[78], chanx_left_in[122]}),
		.sram(mux_2level_tapbuf_size5_20_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_20_sram_inv[0:5]),
		.out(chany_top_out[58]));

	mux_2level_tapbuf_size5 mux_top_track_118 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[80], chanx_left_in[121]}),
		.sram(mux_2level_tapbuf_size5_21_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_21_sram_inv[0:5]),
		.out(chany_top_out[59]));

	mux_2level_tapbuf_size5 mux_top_track_132 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_right_in[89], chanx_left_in[112]}),
		.sram(mux_2level_tapbuf_size5_22_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_22_sram_inv[0:5]),
		.out(chany_top_out[66]));

	mux_2level_tapbuf_size5 mux_top_track_134 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_right_in[90], chanx_left_in[110]}),
		.sram(mux_2level_tapbuf_size5_23_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_23_sram_inv[0:5]),
		.out(chany_top_out[67]));

	mux_2level_tapbuf_size5 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_right_in[92], chanx_left_in[109]}),
		.sram(mux_2level_tapbuf_size5_24_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_24_sram_inv[0:5]),
		.out(chany_top_out[68]));

	mux_2level_tapbuf_size5 mux_top_track_138 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[93], chanx_left_in[108]}),
		.sram(mux_2level_tapbuf_size5_25_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_25_sram_inv[0:5]),
		.out(chany_top_out[69]));

	mux_2level_tapbuf_size5 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_right_in[102], chanx_left_in[98]}),
		.sram(mux_2level_tapbuf_size5_26_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_26_sram_inv[0:5]),
		.out(chany_top_out[76]));

	mux_2level_tapbuf_size5 mux_top_track_154 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_right_in[104], chanx_left_in[97]}),
		.sram(mux_2level_tapbuf_size5_27_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_27_sram_inv[0:5]),
		.out(chany_top_out[77]));

	mux_2level_tapbuf_size5 mux_top_track_156 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_right_in[105], chanx_left_in[96]}),
		.sram(mux_2level_tapbuf_size5_28_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_28_sram_inv[0:5]),
		.out(chany_top_out[78]));

	mux_2level_tapbuf_size5 mux_top_track_158 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[106], chanx_left_in[94]}),
		.sram(mux_2level_tapbuf_size5_29_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_29_sram_inv[0:5]),
		.out(chany_top_out[79]));

	mux_2level_tapbuf_size5 mux_top_track_172 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_right_in[116], chanx_left_in[85]}),
		.sram(mux_2level_tapbuf_size5_30_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_30_sram_inv[0:5]),
		.out(chany_top_out[86]));

	mux_2level_tapbuf_size5 mux_top_track_174 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_right_in[117], chanx_left_in[84]}),
		.sram(mux_2level_tapbuf_size5_31_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_31_sram_inv[0:5]),
		.out(chany_top_out[87]));

	mux_2level_tapbuf_size5 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_right_in[118], chanx_left_in[82]}),
		.sram(mux_2level_tapbuf_size5_32_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_32_sram_inv[0:5]),
		.out(chany_top_out[88]));

	mux_2level_tapbuf_size5 mux_top_track_178 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[120], chanx_left_in[81]}),
		.sram(mux_2level_tapbuf_size5_33_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_33_sram_inv[0:5]),
		.out(chany_top_out[89]));

	mux_2level_tapbuf_size5 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_right_in[129], chanx_left_in[72]}),
		.sram(mux_2level_tapbuf_size5_34_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_34_sram_inv[0:5]),
		.out(chany_top_out[96]));

	mux_2level_tapbuf_size5 mux_top_track_194 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_right_in[130], chanx_left_in[70]}),
		.sram(mux_2level_tapbuf_size5_35_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_35_sram_inv[0:5]),
		.out(chany_top_out[97]));

	mux_2level_tapbuf_size5 mux_top_track_196 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_right_in[132], chanx_left_in[69]}),
		.sram(mux_2level_tapbuf_size5_36_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_36_sram_inv[0:5]),
		.out(chany_top_out[98]));

	mux_2level_tapbuf_size5 mux_top_track_198 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[133], chanx_left_in[68]}),
		.sram(mux_2level_tapbuf_size5_37_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_37_sram_inv[0:5]),
		.out(chany_top_out[99]));

	mux_2level_tapbuf_size5 mux_top_track_212 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_right_in[142], chanx_left_in[58]}),
		.sram(mux_2level_tapbuf_size5_38_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_38_sram_inv[0:5]),
		.out(chany_top_out[106]));

	mux_2level_tapbuf_size5 mux_top_track_214 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_right_in[144], chanx_left_in[57]}),
		.sram(mux_2level_tapbuf_size5_39_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_39_sram_inv[0:5]),
		.out(chany_top_out[107]));

	mux_2level_tapbuf_size5 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_right_in[145], chanx_left_in[56]}),
		.sram(mux_2level_tapbuf_size5_40_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_40_sram_inv[0:5]),
		.out(chany_top_out[108]));

	mux_2level_tapbuf_size5 mux_top_track_218 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[146], chanx_left_in[54]}),
		.sram(mux_2level_tapbuf_size5_41_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_41_sram_inv[0:5]),
		.out(chany_top_out[109]));

	mux_2level_tapbuf_size5 mux_top_track_222 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_31_, chanx_left_in[52]}),
		.sram(mux_2level_tapbuf_size5_42_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_42_sram_inv[0:5]),
		.out(chany_top_out[111]));

	mux_2level_tapbuf_size5 mux_top_track_224 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_32_, chanx_left_in[50]}),
		.sram(mux_2level_tapbuf_size5_43_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_43_sram_inv[0:5]),
		.out(chany_top_out[112]));

	mux_2level_tapbuf_size5 mux_top_track_232 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_left_in[45], chanx_left_in[139]}),
		.sram(mux_2level_tapbuf_size5_44_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_44_sram_inv[0:5]),
		.out(chany_top_out[116]));

	mux_2level_tapbuf_size5 mux_top_track_234 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_left_in[44], chanx_left_in[135]}),
		.sram(mux_2level_tapbuf_size5_45_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_45_sram_inv[0:5]),
		.out(chany_top_out[117]));

	mux_2level_tapbuf_size5 mux_top_track_236 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_left_in[42], chanx_left_in[131]}),
		.sram(mux_2level_tapbuf_size5_46_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_46_sram_inv[0:5]),
		.out(chany_top_out[118]));

	mux_2level_tapbuf_size5 mux_top_track_238 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_left_in[41], chanx_left_in[127]}),
		.sram(mux_2level_tapbuf_size5_47_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_47_sram_inv[0:5]),
		.out(chany_top_out[119]));

	mux_2level_tapbuf_size5 mux_top_track_252 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_left_in[32], chanx_left_in[99]}),
		.sram(mux_2level_tapbuf_size5_48_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_48_sram_inv[0:5]),
		.out(chany_top_out[126]));

	mux_2level_tapbuf_size5 mux_top_track_254 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_left_in[30], chanx_left_in[95]}),
		.sram(mux_2level_tapbuf_size5_49_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_49_sram_inv[0:5]),
		.out(chany_top_out[127]));

	mux_2level_tapbuf_size5 mux_top_track_256 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_left_in[29], chanx_left_in[91]}),
		.sram(mux_2level_tapbuf_size5_50_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_50_sram_inv[0:5]),
		.out(chany_top_out[128]));

	mux_2level_tapbuf_size5 mux_top_track_258 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_left_in[28], chanx_left_in[87]}),
		.sram(mux_2level_tapbuf_size5_51_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_51_sram_inv[0:5]),
		.out(chany_top_out[129]));

	mux_2level_tapbuf_size5 mux_top_track_272 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_left_in[18], chanx_left_in[59]}),
		.sram(mux_2level_tapbuf_size5_52_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_52_sram_inv[0:5]),
		.out(chany_top_out[136]));

	mux_2level_tapbuf_size5 mux_top_track_274 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_left_in[17], chanx_left_in[55]}),
		.sram(mux_2level_tapbuf_size5_53_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_53_sram_inv[0:5]),
		.out(chany_top_out[137]));

	mux_2level_tapbuf_size5 mux_top_track_276 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_left_in[16], chanx_left_in[51]}),
		.sram(mux_2level_tapbuf_size5_54_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_54_sram_inv[0:5]),
		.out(chany_top_out[138]));

	mux_2level_tapbuf_size5 mux_top_track_278 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_left_in[14], chanx_left_in[47]}),
		.sram(mux_2level_tapbuf_size5_55_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_55_sram_inv[0:5]),
		.out(chany_top_out[139]));

	mux_2level_tapbuf_size5 mux_top_track_292 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_26_, chanx_left_in[5], chanx_left_in[19]}),
		.sram(mux_2level_tapbuf_size5_56_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_56_sram_inv[0:5]),
		.out(chany_top_out[146]));

	mux_2level_tapbuf_size5 mux_top_track_294 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_left_in[4], chanx_left_in[15]}),
		.sram(mux_2level_tapbuf_size5_57_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_57_sram_inv[0:5]),
		.out(chany_top_out[147]));

	mux_2level_tapbuf_size5 mux_top_track_296 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_left_in[2], chanx_left_in[11]}),
		.sram(mux_2level_tapbuf_size5_58_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_58_sram_inv[0:5]),
		.out(chany_top_out[148]));

	mux_2level_tapbuf_size5_mem mem_top_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_0_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_14 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_1_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_2_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_3_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_4_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_34 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_5_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_6_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_38 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_7_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_52 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_8_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_54 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_9_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_10_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_11_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_12_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_78 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_13_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_14_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_94 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_15_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_16_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_17_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_18_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_19_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_20_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_20_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_118 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_21_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_21_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_22_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_22_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_134 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_23_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_23_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_24_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_24_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_138 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_25_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_25_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_26_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_26_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_27_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_27_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_28_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_28_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_158 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_29_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_29_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_30_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_30_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_174 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_31_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_31_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_32_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_32_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_178 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_33_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_33_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_34_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_34_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_35_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_35_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_196 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_36_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_36_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_198 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_37_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_37_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_212 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_38_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_38_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_214 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_39_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_39_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_40_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_40_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_218 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_41_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_41_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_222 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_42_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_42_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_43_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_43_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_44_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_44_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_234 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_45_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_45_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_236 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_46_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_46_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_238 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_47_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_47_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_252 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_48_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_48_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_254 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_49_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_49_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_50_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_50_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_258 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_51_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_51_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_80_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_52_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_52_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_274 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_53_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_53_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_276 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_54_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_54_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_278 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_55_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_55_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_292 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_86_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_56_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_56_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_294 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_57_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_57_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_58_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_58_sram_inv[0:5]));

	mux_2level_tapbuf_size4 mux_top_track_74 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_27_, chanx_right_in[50]}),
		.sram(mux_2level_tapbuf_size4_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_0_sram_inv[0:5]),
		.out(chany_top_out[37]));

	mux_2level_tapbuf_size4 mux_top_track_76 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_28_, chanx_right_in[52]}),
		.sram(mux_2level_tapbuf_size4_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_1_sram_inv[0:5]),
		.out(chany_top_out[38]));

	mux_2level_tapbuf_size4_mem mem_top_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_0_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_top_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_1_sram_inv[0:5]));

	mux_2level_tapbuf_size7 mux_top_track_298 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_out_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_out_29_, chanx_right_in[0], chanx_right_in[3], chanx_left_in[1], chanx_left_in[7]}),
		.sram(mux_2level_tapbuf_size7_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_0_sram_inv[0:5]),
		.out(chany_top_out[149]));

	mux_2level_tapbuf_size7 mux_right_track_296 (
		.in({chany_top_in[36], chany_top_in[74], chany_top_in[112], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[49], chanx_left_in[100]}),
		.sram(mux_2level_tapbuf_size7_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_1_sram_inv[0:5]),
		.out(chanx_right_out[148]));

	mux_2level_tapbuf_size7 mux_left_track_65 (
		.in({chany_top_in[30], chany_top_in[68], chany_top_in[106], chany_top_in[144], chanx_right_in[10], chanx_right_in[61], chanx_right_in[112]}),
		.sram(mux_2level_tapbuf_size7_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_2_sram_inv[0:5]),
		.out(chanx_left_out[32]));

	mux_2level_tapbuf_size7 mux_left_track_137 (
		.in({chany_top_in[21], chany_top_in[59], chany_top_in[97], chany_top_in[135], chanx_right_in[22], chanx_right_in[73], chanx_right_in[124]}),
		.sram(mux_2level_tapbuf_size7_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_3_sram_inv[0:5]),
		.out(chanx_left_out[68]));

	mux_2level_tapbuf_size7 mux_left_track_209 (
		.in({chany_top_in[12], chany_top_in[50], chany_top_in[88], chany_top_in[126], chanx_right_in[34], chanx_right_in[85], chanx_right_in[136]}),
		.sram(mux_2level_tapbuf_size7_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_4_sram_inv[0:5]),
		.out(chanx_left_out[104]));

	mux_2level_tapbuf_size7 mux_left_track_281 (
		.in({chany_top_in[3], chany_top_in[41], chany_top_in[79], chany_top_in[117], chanx_right_in[46], chanx_right_in[97], chanx_right_in[148]}),
		.sram(mux_2level_tapbuf_size7_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_5_sram_inv[0:5]),
		.out(chanx_left_out[140]));

	mux_2level_tapbuf_size7 mux_left_track_289 (
		.in({chany_top_in[2], chany_top_in[40], chany_top_in[78], chany_top_in[116], chanx_right_in[48], chanx_right_in[98], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size7_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_6_sram_inv[0:5]),
		.out(chanx_left_out[144]));

	mux_2level_tapbuf_size7 mux_left_track_297 (
		.in({chany_top_in[1], chany_top_in[39], chany_top_in[77], chany_top_in[115], chanx_right_in[49], chanx_right_in[100], left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size7_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_7_sram_inv[0:5]),
		.out(chanx_left_out[148]));

	mux_2level_tapbuf_size7_mem mem_top_track_298 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_0_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_right_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_1_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_2_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_137 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_3_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_209 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_4_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_281 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_5_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_289 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_6_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_297 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_6_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_7_sram_inv[0:5]));

	mux_2level_tapbuf_size9 mux_right_track_0 (
		.in({chany_top_in[37], chany_top_in[75], chany_top_in[113], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[0], chanx_left_in[50], chanx_left_in[101]}),
		.sram(mux_2level_tapbuf_size9_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_0_sram_inv[0:7]),
		.out(chanx_right_out[0]));

	mux_2level_tapbuf_size9 mux_right_track_56 (
		.in({chany_top_in[6], chany_top_in[44], chany_top_in[82], chany_top_in[120], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[9], chanx_left_in[60], chanx_left_in[110]}),
		.sram(mux_2level_tapbuf_size9_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_1_sram_inv[0:7]),
		.out(chanx_right_out[28]));

	mux_2level_tapbuf_size9 mux_right_track_64 (
		.in({chany_top_in[7], chany_top_in[45], chany_top_in[83], chany_top_in[121], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[10], chanx_left_in[61], chanx_left_in[112]}),
		.sram(mux_2level_tapbuf_size9_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_2_sram_inv[0:7]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size9 mux_right_track_128 (
		.in({chany_top_in[15], chany_top_in[53], chany_top_in[91], chany_top_in[129], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[21], chanx_left_in[72], chanx_left_in[122]}),
		.sram(mux_2level_tapbuf_size9_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_3_sram_inv[0:7]),
		.out(chanx_right_out[64]));

	mux_2level_tapbuf_size9 mux_right_track_136 (
		.in({chany_top_in[16], chany_top_in[54], chany_top_in[92], chany_top_in[130], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[22], chanx_left_in[73], chanx_left_in[124]}),
		.sram(mux_2level_tapbuf_size9_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_4_sram_inv[0:7]),
		.out(chanx_right_out[68]));

	mux_2level_tapbuf_size9 mux_right_track_144 (
		.in({chany_top_in[17], chany_top_in[55], chany_top_in[93], chany_top_in[131], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[24], chanx_left_in[74], chanx_left_in[125]}),
		.sram(mux_2level_tapbuf_size9_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_5_sram_inv[0:7]),
		.out(chanx_right_out[72]));

	mux_2level_tapbuf_size9 mux_right_track_152 (
		.in({chany_top_in[18], chany_top_in[56], chany_top_in[94], chany_top_in[132], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[25], chanx_left_in[76], chanx_left_in[126]}),
		.sram(mux_2level_tapbuf_size9_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_6_sram_inv[0:7]),
		.out(chanx_right_out[76]));

	mux_2level_tapbuf_size9 mux_right_track_160 (
		.in({chany_top_in[19], chany_top_in[57], chany_top_in[95], chany_top_in[133], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[26], chanx_left_in[77], chanx_left_in[128]}),
		.sram(mux_2level_tapbuf_size9_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_7_sram_inv[0:7]),
		.out(chanx_right_out[80]));

	mux_2level_tapbuf_size9 mux_right_track_168 (
		.in({chany_top_in[20], chany_top_in[58], chany_top_in[96], chany_top_in[134], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[28], chanx_left_in[78], chanx_left_in[129]}),
		.sram(mux_2level_tapbuf_size9_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_8_sram_inv[0:7]),
		.out(chanx_right_out[84]));

	mux_2level_tapbuf_size9 mux_right_track_176 (
		.in({chany_top_in[21], chany_top_in[59], chany_top_in[97], chany_top_in[135], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[29], chanx_left_in[80], chanx_left_in[130]}),
		.sram(mux_2level_tapbuf_size9_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_9_sram_inv[0:7]),
		.out(chanx_right_out[88]));

	mux_2level_tapbuf_size9 mux_right_track_184 (
		.in({chany_top_in[22], chany_top_in[60], chany_top_in[98], chany_top_in[136], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[30], chanx_left_in[81], chanx_left_in[132]}),
		.sram(mux_2level_tapbuf_size9_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_10_sram_inv[0:7]),
		.out(chanx_right_out[92]));

	mux_2level_tapbuf_size9 mux_right_track_192 (
		.in({chany_top_in[23], chany_top_in[61], chany_top_in[99], chany_top_in[137], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[32], chanx_left_in[82], chanx_left_in[133]}),
		.sram(mux_2level_tapbuf_size9_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_11_sram_inv[0:7]),
		.out(chanx_right_out[96]));

	mux_2level_tapbuf_size9 mux_right_track_200 (
		.in({chany_top_in[24], chany_top_in[62], chany_top_in[100], chany_top_in[138], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[33], chanx_left_in[84], chanx_left_in[134]}),
		.sram(mux_2level_tapbuf_size9_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_12_sram_inv[0:7]),
		.out(chanx_right_out[100]));

	mux_2level_tapbuf_size9 mux_right_track_208 (
		.in({chany_top_in[25], chany_top_in[63], chany_top_in[101], chany_top_in[139], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[34], chanx_left_in[85], chanx_left_in[136]}),
		.sram(mux_2level_tapbuf_size9_13_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_13_sram_inv[0:7]),
		.out(chanx_right_out[104]));

	mux_2level_tapbuf_size9 mux_right_track_216 (
		.in({chany_top_in[26], chany_top_in[64], chany_top_in[102], chany_top_in[140], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[36], chanx_left_in[86], chanx_left_in[137]}),
		.sram(mux_2level_tapbuf_size9_14_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_14_sram_inv[0:7]),
		.out(chanx_right_out[108]));

	mux_2level_tapbuf_size9 mux_right_track_224 (
		.in({chany_top_in[27], chany_top_in[65], chany_top_in[103], chany_top_in[141], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[37], chanx_left_in[88], chanx_left_in[138]}),
		.sram(mux_2level_tapbuf_size9_15_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_15_sram_inv[0:7]),
		.out(chanx_right_out[112]));

	mux_2level_tapbuf_size9 mux_right_track_232 (
		.in({chany_top_in[28], chany_top_in[66], chany_top_in[104], chany_top_in[142], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[38], chanx_left_in[89], chanx_left_in[140]}),
		.sram(mux_2level_tapbuf_size9_16_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_16_sram_inv[0:7]),
		.out(chanx_right_out[116]));

	mux_2level_tapbuf_size9 mux_right_track_240 (
		.in({chany_top_in[29], chany_top_in[67], chany_top_in[105], chany_top_in[143], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[40], chanx_left_in[90], chanx_left_in[141]}),
		.sram(mux_2level_tapbuf_size9_17_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_17_sram_inv[0:7]),
		.out(chanx_right_out[120]));

	mux_2level_tapbuf_size9 mux_right_track_248 (
		.in({chany_top_in[30], chany_top_in[68], chany_top_in[106], chany_top_in[144], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[41], chanx_left_in[92], chanx_left_in[142]}),
		.sram(mux_2level_tapbuf_size9_18_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_18_sram_inv[0:7]),
		.out(chanx_right_out[124]));

	mux_2level_tapbuf_size9 mux_right_track_256 (
		.in({chany_top_in[31], chany_top_in[69], chany_top_in[107], chany_top_in[145], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[42], chanx_left_in[93], chanx_left_in[144]}),
		.sram(mux_2level_tapbuf_size9_19_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_19_sram_inv[0:7]),
		.out(chanx_right_out[128]));

	mux_2level_tapbuf_size9 mux_right_track_264 (
		.in({chany_top_in[32], chany_top_in[70], chany_top_in[108], chany_top_in[146], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[44], chanx_left_in[94], chanx_left_in[145]}),
		.sram(mux_2level_tapbuf_size9_20_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_20_sram_inv[0:7]),
		.out(chanx_right_out[132]));

	mux_2level_tapbuf_size9 mux_right_track_272 (
		.in({chany_top_in[33], chany_top_in[71], chany_top_in[109], chany_top_in[147], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[45], chanx_left_in[96], chanx_left_in[146]}),
		.sram(mux_2level_tapbuf_size9_21_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_21_sram_inv[0:7]),
		.out(chanx_right_out[136]));

	mux_2level_tapbuf_size9 mux_right_track_280 (
		.in({chany_top_in[34], chany_top_in[72], chany_top_in[110], chany_top_in[148], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[46], chanx_left_in[97], chanx_left_in[148]}),
		.sram(mux_2level_tapbuf_size9_22_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_22_sram_inv[0:7]),
		.out(chanx_right_out[140]));

	mux_2level_tapbuf_size9 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[38], chany_top_in[76], chany_top_in[114], chanx_right_in[0], chanx_right_in[50], chanx_right_in[101], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size9_23_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_23_sram_inv[0:7]),
		.out(chanx_left_out[0]));

	mux_2level_tapbuf_size9 mux_left_track_25 (
		.in({chany_top_in[35], chany_top_in[73], chany_top_in[111], chany_top_in[149], chanx_right_in[4], chanx_right_in[54], chanx_right_in[105], left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size9_24_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_24_sram_inv[0:7]),
		.out(chanx_left_out[12]));

	mux_2level_tapbuf_size9 mux_left_track_33 (
		.in({chany_top_in[34], chany_top_in[72], chany_top_in[110], chany_top_in[148], chanx_right_in[5], chanx_right_in[56], chanx_right_in[106], left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size9_25_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_25_sram_inv[0:7]),
		.out(chanx_left_out[16]));

	mux_2level_tapbuf_size9 mux_left_track_41 (
		.in({chany_top_in[33], chany_top_in[71], chany_top_in[109], chany_top_in[147], chanx_right_in[6], chanx_right_in[57], chanx_right_in[108], left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size9_26_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_26_sram_inv[0:7]),
		.out(chanx_left_out[20]));

	mux_2level_tapbuf_size9_mem mem_right_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_0_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_1_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_2_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_3_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_4_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_5_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_6_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_7_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_8_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_9_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_10_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_11_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_12_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_13_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_13_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_14_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_14_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_15_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_15_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_16_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_16_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_17_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_17_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_18_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_18_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_19_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_19_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_20_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_20_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_21_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_21_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_right_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_22_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_22_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_23_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_23_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_24_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_24_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_25_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_25_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_26_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_26_sram_inv[0:7]));

	mux_2level_tapbuf_size10 mux_right_track_8 (
		.in({chany_top_in[0], chany_top_in[38], chany_top_in[76], chany_top_in[114], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[1], chanx_left_in[52], chanx_left_in[102]}),
		.sram(mux_2level_tapbuf_size10_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_0_sram_inv[0:7]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size10 mux_right_track_16 (
		.in({chany_top_in[1], chany_top_in[39], chany_top_in[77], chany_top_in[115], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[2], chanx_left_in[53], chanx_left_in[104]}),
		.sram(mux_2level_tapbuf_size10_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_1_sram_inv[0:7]),
		.out(chanx_right_out[8]));

	mux_2level_tapbuf_size10 mux_right_track_24 (
		.in({chany_top_in[2], chany_top_in[40], chany_top_in[78], chany_top_in[116], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[4], chanx_left_in[54], chanx_left_in[105]}),
		.sram(mux_2level_tapbuf_size10_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_2_sram_inv[0:7]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size10 mux_right_track_32 (
		.in({chany_top_in[3], chany_top_in[41], chany_top_in[79], chany_top_in[117], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[5], chanx_left_in[56], chanx_left_in[106]}),
		.sram(mux_2level_tapbuf_size10_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_3_sram_inv[0:7]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size10 mux_right_track_40 (
		.in({chany_top_in[4], chany_top_in[42], chany_top_in[80], chany_top_in[118], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[6], chanx_left_in[57], chanx_left_in[108]}),
		.sram(mux_2level_tapbuf_size10_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_4_sram_inv[0:7]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size10 mux_right_track_48 (
		.in({chany_top_in[5], chany_top_in[43], chany_top_in[81], chany_top_in[119], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[8], chanx_left_in[58], chanx_left_in[109]}),
		.sram(mux_2level_tapbuf_size10_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_5_sram_inv[0:7]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size10 mux_right_track_72 (
		.in({chany_top_in[8], chany_top_in[46], chany_top_in[84], chany_top_in[122], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[12], chanx_left_in[62], chanx_left_in[113]}),
		.sram(mux_2level_tapbuf_size10_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_6_sram_inv[0:7]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size10 mux_right_track_80 (
		.in({chany_top_in[9], chany_top_in[47], chany_top_in[85], chany_top_in[123], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[13], chanx_left_in[64], chanx_left_in[114]}),
		.sram(mux_2level_tapbuf_size10_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_7_sram_inv[0:7]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size10 mux_right_track_88 (
		.in({chany_top_in[10], chany_top_in[48], chany_top_in[86], chany_top_in[124], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[14], chanx_left_in[65], chanx_left_in[116]}),
		.sram(mux_2level_tapbuf_size10_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_8_sram_inv[0:7]),
		.out(chanx_right_out[44]));

	mux_2level_tapbuf_size10 mux_right_track_96 (
		.in({chany_top_in[11], chany_top_in[49], chany_top_in[87], chany_top_in[125], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[16], chanx_left_in[66], chanx_left_in[117]}),
		.sram(mux_2level_tapbuf_size10_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_9_sram_inv[0:7]),
		.out(chanx_right_out[48]));

	mux_2level_tapbuf_size10 mux_right_track_104 (
		.in({chany_top_in[12], chany_top_in[50], chany_top_in[88], chany_top_in[126], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[17], chanx_left_in[68], chanx_left_in[118]}),
		.sram(mux_2level_tapbuf_size10_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_10_sram_inv[0:7]),
		.out(chanx_right_out[52]));

	mux_2level_tapbuf_size10 mux_right_track_112 (
		.in({chany_top_in[13], chany_top_in[51], chany_top_in[89], chany_top_in[127], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[18], chanx_left_in[69], chanx_left_in[120]}),
		.sram(mux_2level_tapbuf_size10_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_11_sram_inv[0:7]),
		.out(chanx_right_out[56]));

	mux_2level_tapbuf_size10 mux_right_track_120 (
		.in({chany_top_in[14], chany_top_in[52], chany_top_in[90], chany_top_in[128], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[20], chanx_left_in[70], chanx_left_in[121]}),
		.sram(mux_2level_tapbuf_size10_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_12_sram_inv[0:7]),
		.out(chanx_right_out[60]));

	mux_2level_tapbuf_size10_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_0_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_1_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_2_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_3_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_4_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_5_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_6_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_7_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_8_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_9_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_10_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_11_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_right_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_12_sram_inv[0:7]));

endmodule
// ----- END Verilog module for sb_6__0_ -----

//----- Default net type -----
`default_nettype wire



